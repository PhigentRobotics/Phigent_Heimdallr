//=========================
// Engineer:  Wu Di
// Email: 
// Create Date: 
// Module Name: 
// Project Name: 
// Description: 
//=========================

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
GCkj6tr8QkPqP3wKRIO3S0WTEuMTbQhVWmwumMr+VJn2d3caoJVdmDrUzQ2PToGYw2iytq7KcKbQ
ZrlGbzMNiNWCVwY7oXItBjr4qX3dhgnUAVbPB3sLOWmzSsgGqbDeJe5mgUPTfxcwQ1BZenPwvZsy
LrMMxH3rZM1nkGNWh0RRg9AkeL9aU2pfVBtVGsCjoxHThsiPJGzwoZM4EmguvHmSU1UQVnDJggPu
W6+tNkiFY1r/YGIQpSEbFq8xwWtswwjBcbu5tLOUZB0G9QXC+AWH8x6Od90kCCvppZ+vAQaJNcul
3N0HjZ9M0pu/59DFn6nziZ/Oq3XLbbun5Vc22g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="HNcwuMCKZp10e+Tec+d5ecMkvOoxZraTQTUYsHGPmHM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 221760)
`pragma protect data_block
+27Rlo6JYsFWB37cEkrAuzWeNGlFsvTPMKUT6l3LsTXvnXY5D7MUC6f7l5WBlD2f4O/s7beE8ynR
BGNQXD+CdDM9VbF/NqNSFw2Aqz8L768M7vqh8QGY9hMsDH+XJwQeKmLBNkqVbGuyO6wfzpy0lMg3
meDf+tJukOAZYq4BQO6OdVO8v9bZJnqS+iDPCZG/XvkOQj4F+sp8FQ6vrM4jbqzprlqQ+u9QNCnc
LpKe19TJBPUrKcWf024ApFaX9xG0C7ZIu4qcRRb5y5/2vdfTD2zI/7ojrj900buPXVqCLk8BGVbD
wRDAxEXT6YSXPGxjCu3EjbPkWKXylK5aUSGHJtVCel5940gYWBfbxAqhCVnYKpBj3dEMiu72/iwq
P0Ta//Lm85JcFZP0Fbylnbkhpwu1K+92f254xkrahMfCpTAp26BVLkSV4SJjIaYKgdEknOp5Lftd
3Hk6ySN/3/1z1rBZ0Dwn8FlR3xeTay+sYDHUUFj4ZbDrWClUv53edCgb4i0dNFk59AZaqJHLP3tw
zynwtnGbF7Nt1qEjmiBJ7V+wTsEwnOXpSBusEpDXgheL1YvBr+2EMpBq4TKFcKq4iVxnVijxqJ2E
IQENjeesGUZaoBvrSGmvT1It83BpgcEvuDH5KuVHBBFT0bNLjmeQkQUPX0o27EUkP0OMxhTifUsl
It8bkHOJ8PyEi6CgGM/X16y8SDQ8uHmDCcRC3Mn/GiOn9V6MBLsdGONkj2AMaYhvcqVe1C/nQE0w
wGZ+DF/b5ZupFZ1Cjx7vZRvexpostw9pSrtdhAXv/C3rkZ0/Ligg37JAY3izeQyoDIb5R+5PL6Qj
LH7nSS3V9ACHnPeyE0O2I9LwV27Hc5AZe3WgFFOrhcoyGiijkEEILNHH5stbENrvKHu96VeTlgZj
bxNfLCLcSXHVk7UdEkVwb4sjVMnw1MuxRi2JcoPdlWsYDoSc9vwd4Yu39fPhsXU7xOFftkqAvE+h
K0wX7msI8V2A7Ehvq8ykU/EYz3KHMfRExQRqhziyFfjezeXHcjYRq/m8YQD4VTTVRl19IfQCLnIV
hdd9jgDAUP7Ck2jLl/DIswmfl2q7c9XQC24OUOnCJ+r/mElTWfdn/UMzpLgxW5G3gIBKSOot88rn
1tvTjzfIo7hh4aUzlhh1PsH/iTIFLgUkMGNADjxvPyOGRYyuqsTu+A7xPmuDmBqQzCGWnpitSb/7
P2DZrGwR2nQViqkZENidklSS1n2jFkj4zzm3JOGQgL9es1wvWt1WfGf3azH9gjdo/ajhWnsSPq8C
gwJLcMXeeChiMPp28mdtGg8Np7eS5QhSYOJ3u9yIvxWMJj9N3mmGYAwDJASSThL1YK8yr5jGPQUi
6uThEtI9fXDEh0fixawptNNE3pzGBDZA4/2wMPNGUNR8RQcWrFxTg0RhM7yLQtOrFUX04b5FyoQR
5qVMdh9bFxoCwy3F9E7fYm+3xB4cTGNv8m26ZDQUNbbLQaeGDujksQVD7g+xLSjbLHwneDm+7B1X
58NxgesuFxWrDrdio6w7aWpckrjxSXEdzePjrUkkE87t2DamDFKshK8Ai0tAHe0g6YCv0t5B/Af3
65Gr0VC3z3xWqwgNGAZnx/+tFHq1XmdKTe+FRTPWrxr6KKZ4URKdv7j5F4+UlEn7HP3LJTufQ+vH
n5V250TiB73dBKSZCZCxbR/QEKhm8BXVQEl2RImL+1HGnSCrjROsDgS7mc0vMaUmJpOtZq2sh3LU
vYMyw4A1a6OyBUI2NO0ff1HLDm3UkO3XTzebJQ2L5XpfG5LpoKQfFa4v8kRbbaXW/KeN4Y9ef1e1
L975kFLSMuvafx3m7GoTuNZdrkaLHjKsXKw1OOGAuJrZ+JucWUGpzBJOAtcrBJKYO1wkG5bMMRFY
cIE3ylBxUviqf75v1VYwwcfo8BaIh3NxfVOtPLWw9zNTMqCkpmV4+1YvP4h7vQvkEzfaWEA8zCIo
hmYiZwYKoE6BghfRFa/lxR5RdjaGYf8ZZ+pQQA4fmb82/32x7dWPBWZUf3Eu4lDFSDh8aUCRdHlz
bAzAtLLLoyn6EM/nO02Gjd5GSH9Nqkytx/fRNqtqKtKDZmVdlUjoj3deAPl8mof8fX//dYTBgfNg
R15n10IYK6RRM7/nzLYJizQWPkoYEfWsc++DNG1MkG1+nxtQ5fvvagtS4vhKo+3TKVgtjtfQwxj3
IMjJjARaaN+SgkXYZ9o+LP641vXXnDSRyVG2jqr0TYbGmnaJ3ImBp5o79YuTTAxpRDSiOfaa0ZGn
ZdQYe1ZFbh2pxg5LVeojfj+3dW2WVZluJcZshk+WUgHsaMPev7SDfjz9ciVvGypZjSgR9X3mdiz4
Fq0FoyxF5ts2Q6YtNDURKcAJvRqfEDxuED8fP/SKTTB/poiPTeLtyygvkXJTaZ+Tc077XJuKGnxw
iDRZCJEvsTlJO81++X4G5EE5YR9fjFmodD3/Y922V9DRaVkAWIY3YMOO9O/HzVGfQTEU6vaNDAWm
rhigkuMzyALtItsbRxn36E4utkGlojUjrChNpeCZbwzPQjEtMrJBwZay8BpSSSQUfk0XxIBjWAoh
jcEnSYbNtG6ie1AxzJVVkzyz5FQsXnzJYI88kGem9V397srET+AZnXTnsT0iBowI7Copl0epElDe
40YFsQzuAMVC9jd4x02iCFxULXpgPCOAWNXbh/IXWw70Jjmv9krIOwGkgJCbnj7ohXqx58mqjBW8
hDQRk1FWjOXCgNVBWMgS2W9Jar+drXyBs7ZaU/IWhE2HyUplBbpkvc/dWcpu3H9neKnl/kRbRuw5
41LHmmoXo3s4l05aqMfP0gezFU11W59F9F98SeIOkpCHQNnKqsVdrLRVpvN3IbOfFdiRGZcwgG36
mCky7nsSBVYqdzkTfBs0qe1nRDumUMJAhkQZlx2RMz26iToWqKwXsP4Aqr+nQtmfHsjZRZh2Qc9w
/Q5te+5+myPy8L4/csOjFu9xn0ytU3HQlv/YbFEtIEkvAZNwep/ioiset80WtFJcLs3wcgPsR51X
CrLdfCwsAERxl5qTgYBYpdUCA+pwYTeYkMp+ruopGuOe5EubNGp7NuaA0drtAsp6G9xxlRAF5R9E
ER+E7YQwoM78P+ok2Hi1E6bIa1fy97vNCXdekJnUzNf1y748t16M6PZCC3KwN1WUQSbVvDDtyniL
O2JX8e8IV4C5SpcvIDpTe4ld1fxKSkp2vEhd7TKNuyZzZxSPQpdW3yCGnAWUjQXwRAGPADUwQzqL
Ep+3ijaSFp+bfS7N2o24nmREstJvijnZ38AjoLsdsVtcua5YONorWOKfT7vIlGSNiOjANysvMohC
rfCP+i3COHA2al2uuPgI1WorwSvdi3T9LexbaEUZ+yR3j0qUITf7O3g9KkadjOkLPTjFJVckqoQC
UrDtMZh8zUcNFVJuS1Xx5z6CiyTV1jhj6np4/W6Y+OhIC0w0NaXZkwzIZAOkcsFpol5daMbChLs5
jPRhau0l0uIZRrgMyCUAkMGc/YYoPQ/58VAys+KKykHocEw66oiEMDBjvzjU2cUYdqjtG5vOF/g0
KZNAyiyAavy2DJgWc9ChoNpgiTG83SY/PEB/ZBWd62Yiiyv8OWQo8vGsW38LO07mOjD5o+F3nV0A
egr74q6Y97v/klYJ8LxTSP1nObxCv39jdfMtnEnjYmnITqTOBLPnwc6a58DyygfMK/wKdVlV/k4H
WqgjGEpmJfvcRt5ya69fPrpQSx35wZUxZIYqeKR8sun3QEjWvzp+8pyT3PDLcmRGT6h7L9rUvCKp
l35XqW4N+WhkGlDQaBI//2lqRZLAQ15pKmTi+ra0H3VmzBbflzLcD5TBhGZyQlcqsRTMRHbv11bU
LZgikn15F/GzV7Izr0scuH2eEf8Ytpdq2wrX/Uk3CWdsAQvQrlzmntsVvqBGjTaL8uoiOo9TyvLZ
SUuJYlE0sqMFP7KyqO6HVnzJDyouhWJPiVGf03NxIkKdgpTPb/ZsMyUADHT3+iwl5CfHj9N2muqx
YBP+0uMEJQ/D7CAND5+X196k+o75o5Wg+EkMv4l+10k18viJhmPlinzoKggfZaIxWhV+dxXslKjY
X+eUD93AMv+kLfy6oKEWb1kxHHpH7boYVzsvQI3ZgYXqFdEhJiFmkPfzWOjjXzkL7lmcThp6/ska
ZSx9n/cV5+EzVGnqSoiPLUww9zQMxkIEifFXtIZmCiWG0UmUsVlYCsarNJ//pNc7mgw9pgUejmUE
1MYO2PnA83jgP0aTLGzgKTchQgjz+Fc5Yq/2wcfbdgoX9/OMICjxiPuOzuIWuPr8zvWaeUOSWJAM
siRhcqkj+uAJmE/QulAGqF0oIB9y98Zbo13UI1+xbBGoOMCM+joGvnBo9FnJ6Mwtn9FywruDJWQv
wVixQTWVaEJ2IxQMru39FU356pBiazOzFdAFSjgd4KNy7LtmZv8HxLjTGR9ylqLjYQgG0EJYmeFG
llvglJDQh5khdGu4n9KbqfPy+etXvnsa/i1QXCr/Vlt7/1TEV2VS5EDl1BURt0b3rlspfmKSa7Qf
AwbRLzPWX5pQ8tSAJeykFbAkdHrdHWcN+WGQkDEaeeqUzrYQ2CDSD1TULD1igEY3PJM/Dd6HTexr
oNxRx6nbOBNTotPRNYTjfC2mHKoR7g4+h4c+P7nLfWp6mJITWtMQB2dLU81qZUCu/vuc9/tzGTwM
rbL55ArOT4oc7MCI6wKwZEu5AVZe45bf9LqtVF1dCAoV/w5jYctqTiOnl1DoDcWeKQER/bm1Epsm
p75M/GW8+QReokDGmMnvTTPcE1QEk46CJIaBcXYJT14sGUOIztOIFCS8dIJqFftUvF6jTHtMQvFT
16kyW/jjcZSTINd309pZkLAXaTq1J330qRArfbzW8aaeN6UnCCLR2GauYwihab+kJLhAlauYucQT
voSy2VX1cS1bI5t7PkMKdN/crfzSqnEZpwdoxGrDaBkoLeX4SvIsn/LHEqlovNzbCwd1zco4OCNi
bEQDT9ZOQCj4C1q6jUn7fAMdRLqQNpbSh+LZRx8pg9X9DI0RG1OuAeQoJabrWeVjv5VHGnyX8siZ
4SYcT/Q2DNyRs+5E4JDVzehIIpsGCtMFsqp9IzrujogF/J3P2v30A2EX5+k50nA3BFtz4OjcHWrc
Vw6LSNH4K3ZFP2GobSD1skzxeBycQmso8CTXqx+rg/szBmgd08XxpPV2U0ZwD5qnn5CphxEGv2+I
eBPGUFsrXZUp2megNtLcGpyhfP/jTuWrt2NuylJ3+fsw2D2+Xurwv3FpQIdZK5/VK1SgUATGLjFw
WiEZ/QXoBA2xaYf7wKbu3xgZa3/iU/RnJVGl6DW0tC/X+1AM1HrIjXWNPaGi+2R/xLLpXiPl+/06
/mAPyjtMrydSEUjrtAWSddmveHb8tPukX8pfBgzOfomcViY6q6/FeGww+TMzIly4G5+tbgG9RQFF
22ldf2HXXrmT2sqFtHscbTU67K1PHPIFzinyC/zNNQRRuKijhi2nGQTYoMqAAFgxbV6etqb1k9zw
HQATc1Ed1j64f6glY78XHcD2KuXEEI8bQ7gawP+aupvdGNAqUpTFi3QOIxzbxiFHpzp8gFs42kQr
6eq5xdaWyKnL+nBnP4BX2o8NNgn9vVDgOoXXA3ZKcklTjXJb49IayIU6TXXaic2XMQdx4mSjeb6z
3x0vJKIVNFCROzAY3VoG+52fmd3DMO18MV0KIQJ+dvZwhBT+IkNUBY2Hb6koxi0kBEnoEhFMh9a7
XDg/rfijA8kplakeYkuvEcmcGXb71a8ptGTOShJERC9tkUG1fij2/ua5S6UWlUiazDKscPmMCR5D
LGa7deymZ2NFPoQXRyIjOM1xXPc1r2H6/IP3mOYH6AmXEbHESEWnwopoy+9a796qqYMlAkPdOSft
04JcExCwv0t+cFbOf86XJ80weSAS0KtB4TUjMlaESLZ4vaw82YFprh77qGls3TX/AhtoNFWccm6x
PEvXcYjDO0enp0feGEMWBbxqikcRSyiZ5AjjOMte1LvesU+DMR0k2C+tDx1JwIMMYA9+RLlW6Snz
lyEQHtivlodYEpyppqq0Xz1vrv+JSYBaJIDKpLXQNoPKmpkDV8iFmsvfdcfACHXacJSI3ZiQIFdE
6/BrehZddDSCcOmnhKJte7z48ZEuK7MWV8WPNUOKnTbeUzydDJW2FfQzyZVDCzCGJGx0eZXIp9XR
txaI9BUcOW8TIV5xS6HnYsE9DDQS/2LFV6SIH2Dsur3ELF7LucPGwICGDV2IxdV4RyjwAak/edHF
SnQup1R/adlCRwAR1pC0a47Jk6TUQTRUnwYEktmIw6mGHAts5O3YkVD0jRl9U7+tPH8/djWbvxGY
U+2lcPPOeImkL8wUPhU+4UKoKUc0//F1hgz5KFRH08g9JUXul7iWF5QZtxHOJCh1y1yqTN6sdwKq
ROSfIw6ZBUBjrCld5vEcF1k2x+hLAfBbgTPCuiI6+ltX5mLOM5DH8i0BONFQozx3tTOirJ8JBLNR
PYHSo6ft/AgnOlma0+S2AN0WTKIJoWweIHXMjtTHdH2NNjjltUMvS1z+dg6cRHsIE1vpHLFlfuqb
DSt0qEUIjDVccBkbZQ912a+WgNV4+2ns2dOZnKMi0y+wXvCaxDXxlr9MTQPr5+iJv/IfgviEyJD6
U8SyFuMpxig8KkHkf6AOQBa3x8LlBHdsI5tuzEvLNwRmGFZdO/Nrzhyqo22N1zfW9fxpR4WpuCmE
Lr/XwbUTZ3wDlpHQjr85f4vZpTbC/fMopMpTM0OUoAHME3FGKZWrL6GGRmKnFzQnQpOhGWJ/owc6
871NGc48DDC1GF55EVhhw94MXF+vIuSbVCOzSgBI+Q1jOjU+zBdyFc+sv52gPvqogQA41v9GjfZX
Upr9XyKrM1StcbSxYE2nffayKk84vTAP28QmdKFa5NfoU5q+JfuWzTQkeYET75k+ecPjFu2C+pEi
iwbNpm6/vdGAc948JiuNatwz9bJsx4Tc6yNtzfXjy7wUorlUnTH8uEuNoD2ddkc4H/uRrHH0M//s
NVzHx9pNUPt4iefRy26wxExa7INwkc7GhzLARKs6d8sTR8nZINWBepT7XWvLJ9fGAh4g7g5Cublz
sush1hA/KWKJ7ytq3ToaQcjvXCP08hIHmHpM+NGZr/lavj5SU4HbJNRGbPChF3cple35K76mWvnS
osa/GpzKVre2jyADD8uWwTE1twB7VIOFuGsd6Dg742Zpv8wp+SPSwvEofQy+VPF+toRHECzHCw8d
LqHqRMk+2+0LmMbOEcwFF3zoo8OfbHs+g3bSFxXA6QfvBoucwEtO3ibVARpY3Pz+MIjbotGthf4D
Fxsum8u7eeuVSeK6dP2JInNihmKSf9hfQw6rCDujze/4/wrhe5mQ55ke3PzhUdNaHkJQQ1z5zERB
QTOrdqMSIGoMYEuRwNMBWJGkx2JJeP6jwQCy6F4M0/6BD51qU84qfgcb6zcog7/rrOVVUvH06zGB
XavEUzFlEeXjKaluRB4ltojP1yz7PCV5A0r94YJFIegN5/yGnqp10Yaf7y1h7XjpD3gD4DhI3ka3
gm1O6t4PB3HC6RXJDflx6gMlxZljg3L/8NATXXQQQ05Ejjaca588VxAM3/O/g/CnJO9X10pZgJne
TIPNpUsQYGwhz8qcBHhkIvLF9X9AHHVE9DUyHw2Hyb3LhbWzgFRZtCdyAiTQq6o9wANXx6z5yXd/
3xn9mJmIgN1JGmQnrGQGLZifX5GtiJOG8s0RehUZuBoh8to6p08EGtD7jjFiIPzicCN2GuOW0e81
JW2h/uReEqAVeOvFZWneWLdmm8LHOUwK7E/xu6V/tejW+KOVQys0RaodQLpYkNwVZ5dsh5KAq1NB
O3HqEGnr55Z904DTu2pfXmoC1Dga/wrD512bjW0TpMwJps0H/x03MqiOEqXREZ9Xb+bhR0rqdd3A
Go5yme/RAl0UttcUlSwMZoz8MVg29eNiXn12rPNvW8Cj8yCPmIpAoSAWV17ovZBqm1i6g/sWRTU0
v8NCCv1LrmMkev37k/Tgy2yF08cnn2QFbel80D5ju6CNFykp8R7wjCvTJJahwuCZJMYDJnsOroz8
tsdeQYKBJTgY+RveSjl67tZmh5xlTYijB8JrdbjZt9hGfA8300Q2Ras6N8DqbjDSxM9vVHa2Za3/
Rtd9I4lavD6Sim2ozx+VmzFl7hkRKmrCO4NSjYJyMfO4SsaEf+lrFRFbLYbleSZ3mgn73gcm90Si
aWOo4E32TNXAk0dw1Lqdsyp5bXAix4W1elxbJVuezlM+6v2jZGREH63iKrnOVkkPJAy+jXo7nFcA
6Ly+Qz7poLKyyqvCCb3UxtYSPk8DIFLZwelaGMIEA2SBHbFQGzTzr65DCDptb9W1UR9H17UbNbiD
IsaRHb6bYEMR84SoqtnDj+Z/wPcfZUt5WUXU5WZGYYkGQQEnDIuYjhZtrBwZU/qkquQKQGSn2b9K
tQjEhsJF9Fa+XRUz38A9IVhdXStV4eKA8gPcc3iLR0IVWw6yLqC0qMWaeQw4ORIoF3Rh12ka4Jv/
35VdU/sP9kxkqCc9iGf8GJCmkOvhEaDrsGQCQevRub3+Pchc7NV63EZ4EObK5gKYVpv59102tXCJ
9vMsxVMkU0bGwa3wl+Aaa3Oz47jkntBrCbx3SUGceMJ0Oqv713vLClK1XLKYhYhHRWCTCCNNNalZ
xvOjsKDwPhWwiHeoevPKogLgFRbbRF0UKV1AtKp5qZdRAdRxQIMk8QB+ZqDp5820WLQDcXaALvSE
YmkKZi/wNI/7I68DYuPV86eLkqKXlAenU6yyNW22sB1MDAk8jNQd6bmuSmZyNOmjkIRMmyQNR2/f
JWjMmTahBB8ctJIfM9OSeORJyNRDt/mTvdMQJ5JOKzrgWE5pS/M/aOnIrA4TcMn1Aafw+gs+0buD
9DwSoLkluhBbtNds4a/+quMf+RN6d0dSK9mTY8nX1kK4v46P9xM2Ehmh0x1B2LIQ74OuXuDyRHSQ
vEkGy2lpIVwyggt+kjzev5iyu+KioVMByBb0lLPgz1TE8WlCPYW2jFaV2RgTddiCviGfvGg6zkVT
kV6/+WmgAwiEU0hW0pkxfaiXnzae12dYX2BOmLMItncQwOzk0UP3KqpgvkqOekO9H1XyfEEUWyAJ
9I9jozWoncd1fGTPgJ9pBs7TZQUEyJ8Fl79VERt1aieZD74XNhZ2MtUO7xZIqWQoTFM1teJhuync
fswCoskS3Mjr+7nmCyhEBX8bQZZHv11XUb5DeDRAhpGYy2Pn2uxoNH+MFwhHB+b0oe77kD6FrObk
zjdfzpqWyXMfLRiBfXaj8XEmAHEa48+v8/68o5Pime2nAzdYI+4992UKr68BTCG3bD2WpjeLr80u
YI/ni6vK4+6LEn1Ux2Zr50875F1Q8qjFfSQovepTyaDef/3VlPAR4ILni0TK/4pDsnC74cBmc89t
E2RVDY+PLNIGRtW0N+hBMs4tfWUSBrdS1KFSHYoAss+7cFIr+b/xMDxbL1GKyFnlyx+wTQsojfnc
11fPDSXfNM47rjVNoq6AIJsVJoJiDjLCBO7MG3ggFpZibY185pImSXF0EObrTiypNkQeJ8scyMmv
Apxrf36MKO55/cCmCQvsQOUKwtBvpRNvJoy8axh+OhVKKnyj2kKxqJ0ckwgy2tRelFrn3IC4Czt9
+8kqA3HYME3lYmVtEIquewmG3gTb24/lGP4btpkUFkNCXfb32AoQz7chgTZN0YFyARZTKBQsWe51
MgZiPxbRKhJ0uaZAr1V4WNYv0wXtH5KBXPzpCSkCZ0YG23ofSf/ouj6R4wnscBTtMPwsT2FfWiPL
qw/gNSSHjH7DhIttAyIyUCd7g1nVLBWVyJkdc/NJPl90rcNWGxBIGBqXSyxMOxcHa3UXn39Zd8Ck
L/Z2pfUH3DjO+W9sX5UqQJpUjBYWlbNwaMmQgdTojv4wWRzakSg2VfItzUX0P1f2ZXGQBhL+3Ely
LO8tM4aKoT1NBH6vtx+EOLos6kJfomsI68bPXwe+kyIxZH6TprFRKqFerbrUL1n48/iKgPJdMGlm
FTsQMBW9gzkxwxA2YgqQJT1Ck67GhHFo0POsPtjL9Dhcoo9E+5Zf2ENapIFQeu9b+PlzPBXLBH/U
ziS5rKk4+kq7oMCNGKC2aAqNfHEkK16rpcVgjz1rm14Vx9qj6IB0qqyxEETkt42d7T5X8P5xdbIK
8GDAZ1sAI0O7p11vLfU2y7/3ynlMx3+Tt59Iksyk1axgzcXQ7j1gaaHVFvjEzhWGvbrolCHPbUDa
NlpAMKUZbFqHwD4wQxjzcoRL+8UfWtZAT8/Q//Wf6YyR9R8ieQi1Q4qJaXNymppbeH2Gw+HqqRhP
T81jaAKQul4ho43id05lIhfs1ltnzASJO4uh2vLd7mGv+rWO8FvesaX9rGMTe1AZSXWk7SlwS++5
g005D+R+Xljkx4SCsXHDpbRtw3R0jQ0aDFXY1DBSy5Qt/otFK757IYw/9FCmb2peeHLCo95uoNUT
ytM1Z4fbrlHJ/DJeQosl0FqcLOhOJWd9fbiVeB5UUe4tWG0e1UfuZ6HReFsGsNzX4ms1v/Drf/Oq
ckl+970Kgzj9FruxX1RZqQx/iNSvOrk7g5mwGqmxPXU76ua+HTEgR5X7UOGXx6uy0P93WtVP/nOf
6a0Mv/xjs1mC4fAVyy+JrsRAzGzeSJoAjmBjDgkmeCrG0N4wmz/6dymN/sOo6DmcSk98jlaNaKio
NJWOngk/g24wAhr/Wc1BqM7eyL34ZdTIXIbaZpkjOuT3rYc+DNU0VQ7UC0z9KMICHu55j/aQnlHV
+H6+QTWSafllqGi4TdIE3XhJWXhC7bJgDrM4N08+ZvlDTLKdg38h1znJpAOW90yUPlKcDWp97DJS
ROU7roBbgxDWH7aiJTkmrXPli9ivep3BcXGDM7JkOAPAVmYXPbH+fdQYfTHRm23E4rOD4rHtemLQ
Lk1Z1LafFYsLujn53zN28GAEe8UbtQDwmsdHRvpHCxNVuJ5eap1In2D3ngUeHoLMMvxpy3TOmroz
zL2Z8rvTmV1bdj+1X/yRrc+g03376e+JIKVhW0+kfXCuk1XNI4ak/v25xmFdeGnZTXzf/3+86M9S
YidgOcRng6T2C9A7C3WnFg7pRkCNMi0hPtY1HE+sKhZEuumeSAu2GiEi4/5A1fUl/QqiFKepMcWm
eyEepFVdE5i0e5BYDyl4eTwy0Jj+UmNUzQHv/NCzi1IckzgCP46C6r3H82u1Wxh7ez8kLuDy0adV
GmNAcpoT1g3w0wB6DxOM0X2SEWLZQLtdfU4H5bDLlpevh2gvSgWnHieNN7uuHMgMuY8rlHaaDaxV
XZaRUgGJu4/dY+t8Gz0YPw4R4mBluTC+2DeBnf74BzFOvj3RB131VXIkGzpAv0Z54v/3s1UdvRmy
R2+vNyOPTQTa+bsNcjLlGEQNaHIVoe6PubIuxftRUNoc2VWVM1Qd1+3NSr2CmbczdxV4utxByK56
Sjj6txHysgCjVVotFVlkAB1ZymsFjdjPag2zspYgLIujNjjB8i0MVKL1nAIMCnft4yrkvGuJkKLK
0PavJy2FhtTky6O7UkIFrpf3VTyomRTpcbI+6t3gWGGLmsecpOlpmftH9G4YISx3DTnypTnQWzcY
9EvMVVQGy2lPWN4bZsB8Sh8OLCNFWUD8tm3pxAU4FvuNsHfQRwAZg9RkmQkQMuWRVdhD5M5n4EZs
DOldWuiNViDp3M/8DzKbKHJe0jCuZhuWX4bCu6ijiTP4PJa3DzXLejWJJHpskDLIY/j1Xh1nAExU
yBaOrUI7YU3WB5cyPRgOk+EsfpGf4f4yAfoS7s491Dk4I/DDs0BAbnA994b6HDJpCM5DXsA4Uzv4
i9gFThLmsnDQXzt443lMkxztJQzLY1orLyBW+NFW/k6s4mkL2I967TiXlD5PwV5DVJZxn9JowsOU
TPMTbUHWxH24YqYS1dOVLP1ZuWz3aY3fMTYYJMylszMT9I1TKkJiDnkAHHn5ACrs2viQHNFRSB2U
+I7fascNmszWX8xASNdOmp/zB/EQqaBp5CU0jEIdpw9BWDbEvvreNG3byHh7NPDOp7MvA7DnSdW5
5IyvpokH02WV0jfEmuaVhrQCGRaQECJr3Bg0mjdpSePD8C3gsaz87gc609Z5whIzD9H5hNymCBLA
XtklP6BOfmLvA+xFECccgjiBZ0ACCKIxfAkD+d3pQ3BUBFm28Qq6KW35i246K6B88zl+V/SK7Yxh
cjRRA8zgeNqM+HRj2U56DUMI4n7LK2xUbJM6m2OU7d76MOmNqNuZ73VUYEVm6yYnWiyEJS65AJ23
c1If6HFp9toCL6sl/y8ose+btMPcJCeNv4xpLwQUrUQ3wxQs0NAD1ASIZI1fVXppf29lW28xviTw
0NBarZrtwKSY4hnTAK4SCL2CrYi/peTgDJCcXQFS/vaIeUhUxh2UYrZj7EG30NbUbEi/ggIYqk4x
MeN+tiANFNoD7+6rks/r2nqbd8yzMxX9fI7LRx1jKAdta+aGT9iV3yHoItFPBaceYNfmCMEtClic
2PWSaPQExTAhHbjNgcAw7iKRm2+JibUGCU9QiSp8okgPwqhW2hcSHkvs5zbll/FVt1RfrwPiDM0x
fDpyUQVoumSXcVaq++B1dJhUkvDp4yhpxCTNdQD5uoHgGwCX9zp568tVHnrjyKwgtFZwVrqHJb0j
lCk+6l810HoDvaQ0Q5gXxAokIfENgUJHDCVxhDYq0z2EzHmbLUEuwcXP6Ks3rm8FNr2mDf2ueCzD
eyiMrOJs06tBuRaxFc8ty+/8ehiSOs2C1xCwa2RR1wN3f6MpOYgapD9Pz5Jgt6MGmbiYE0myl9MA
escPhlK7ktLCVrnHZHPmC0qLERiU0T11XyRxacmz7a6fhCOGSDRxBX8usIljRcydLUZMEGaVSUQt
kGIKs9kLZhmLVaL2jEGKSsoOe9WIRgmxNEAdtUI9M7TS2Z7nXMWAx8+dwOWNreIQj1mt1O00EN1q
jE8XGtwBq/Vbzb0I+Q3WTOdyoOt0FAH4q3mwE+s+OhVfIAlRnjk4IiacfEYDynxsD4Y9uj6AaZ75
bYz4fn2YGtUCVd1n4klaWkaJQAt0DR3cXQQXISS6S8z8LwBIN/kXESox+ln5+OCfYFGzch2ejpbg
t1rkvX8hr+g+7uwFeNjWt+I7irj9YG2VFlBlYPzKFmHtnDQ3ueeGMRdIw8cj1FoACY8zotS2W/wB
zKmNwOSBmis03nnefuxgSqXBvytMdTqgak+pan0s94sPu/z992G6fr3T4ZZc5MDXoA0CkgIFIVGy
pHH6Zen2R6ewvJKfMLQVDdFvP1cgxHaqGOHpCJIQgTX7FNLOaF7smkUeoiw3Ywz56SJ8CGXTCroX
NS1Sz1qqMhJzEvnU2SUqp99CSv4GXf4Zi4QOvQTEfuRErapqG+IYNk2zPWpc9nJDUnNWfM3DF5YA
vEdlf5pisX4XHtBODWHEQLoAAzhoTO0QFdFfIfoXhqnjk9dA2Hq46Xq+8rNuV+OrrVevt9ZVANec
/kV2kNf59rjIRPqHHM/pmsnoeGeAv3p97XHmd1W+zHeht419IQn85ihLbZCRiNnmRPiHafQVzuPP
UAUTgU1fat2M6NtVnf0YnbDbyMDiQosHDHXC2/1vW8uDpZ0NBywV3bJMcfn2TzxZLJ/+nE04FNav
xKUu8rS+iQcEGp20tYPLXdHP9M672cw0Zuw0XZFLIoYMICZuWWixNaWes6NVt9k1AH3UbIS/KFdq
U0sFWQTSONYi5o2jxegivkrb5ItMVhTJC1gdESWUTf925+4NUxqOFJZ8GscS/W5S3pYFwMOHrXSK
rwdylOrZhFFy5r6GOMuoGk4XF7It5niRXkJZpsllRSlfBzGi3knFSSCupgzCVQhGuqM5TexuoqbD
IyfIwjFKTAq5V34aQMI2YDlhdD0RA/AotoTc4IKDqO5c8ghJWU7FZcUXn0+PN6tfTeEi1R1iv8k0
SiG6xOIH4frzUsHqTteI/OeGFulSsZggw9WMrkQrkpGAnrYxyGczqpIuBhR8r+CcCKNX0dBZvNol
VWxACu3msnIzi3jK4JeCpg60GaIFk1xmhRdmnFWmRL7g+Hkn++wyiRTDZvW3pyY0dcWymuheRGiz
hoP7j1MT5HlzyWNGj3oNG9sGBgyw/oLD2gijVGABZTmtcL3cIMvljF5lqTVcM5xwAJ/oeErt7XHu
8TrShOtnvKUGqg5Yt0EGq8zRgbB9EuVXtbIvkOXCv244hzsKHVOXJAXMiXsxks/ztfJ49rR2txGZ
BOH28LKyl+fv8G0cSfCxPH0yHpvoZ21PSwyXFNy2P9nfv6W/nOF7oayJBKGwBAMe8T4zce1tiGgd
eqek5c+YvAfzxj7E1eS2Do48PJ06MJYnvil74hg3g8jwBCRBZU5P0E9dwCbFBC98Ol039w9k5U9j
Dads2luuxyMUCrhJrqmNpzp6walAuDumOzkewGmaGwFuzf75hAOhsIiexwSdcXETN4j+R1Zqg4pb
rGyd7mpN7uZaRlpSMynvfmZ1voRCErJqYilxUZMuIKxKSA3yBEIVnL2uV4888pOG/aaZXpornncC
ch34s7nxiz/hgRrS4PLUot/+3CxzyboCWZKJJgu6Fe8NWhmrLVaWgyvQvwZKGmupZyFp9bACzUcC
mH3SekK6S2VM1RNU35gNeWGBx8rZmG9YIr6hcCRwpeYoHgBJMt+anZpacIVT+u4qjY7BO5AlzB+j
4sbA6ZoDZnbqY+LuyFnQUT5mDpWtQC8L6uLV3K7LytzAEv0bG2WMAAvP1ZLk/653CcRpMzLf25Z7
NRNepvJb96NQP5FcnGRQlogViOv51uzvdbaV/clIcVbKZUYfegeo0z1KR9k9DlkBRl04v1+yTkns
Zi8ShYwhYQvmhdWTvyw5ITIbotqMEJ32m6DUTqX1Dq0z8H3Xm3FLYn5rBgdOOfyY7EBd2E/1zYqA
mVqlVMBIZWUgkkxPny5Ti0T8HkHEaanzbXtHa0p74xhL09AvpEgcn207rkX74OvXRdRCvIu8Y8b6
sOKRtAD9QfCJdiLqlXOpiLZsMEofcj/t8MaLaOWE0+sMqwVEMGmryLBSn50hYpwKT3Eg4LxPHOga
3v4GTsiCbg8YmQ4E9xIPgciyy1LjgY7EAkU/Rp9Lia/1uf6IkDUZ+Gcv2v0I1J5s+WxTsy1qZTrP
7jr1+kcwdMI68MNxpVFiyUmiUoWO7mS/0L4649k0qAci+vTLDtwNM11ttDOdl4WOgTP9Ur2C7RqG
w02EAmwu4scFrh3oLypbjFkL8tblzVm/bLvjGiay2tPsUlAyIcHEPxolZHTaPhBooNielB4xih+F
v3WRjk3CrFz0s1qDIUqnCC1M6uJDMqJNTfcTaiKXaF6x9IPT6L/1WLqMMlUgeF9WAZ9733Bj+7X4
wNLiblYiqANZeyRn6IpGZ+P+3EI2MkwqQICHgVq6gbsUABAnNCSPZjioi3FyYdT2I3dhgCACrnEO
0NGSQsfg2ak/upueI+6fODjQQ4B7OKqGmOlNcIN/L48yuhfRu1Kcgwnf3n6qOVXJTK7sZWzSfYsV
qvCAobQwu201JRa0syH7vsSlb+VmB+aXv2NRhCaPLdulEkLZW+M/pm95nUlZ4iMyXeOclgbCtC0J
perCmJ/bPETzDX+7xrUjCbd597HA26lgIPI6hh9H5QwLudp2/H6NyjQIMxMNRTlODwMHCvaWZScZ
I09w2NbKWD8n/H17Kq6TA8s0o84n/4rUvfPc51nTnBPIhjy+44MXav4JeVbAJ50/FhMVvLQHAhqk
czhSs8IGw+wPbcU1ne9fjNYBSXYM7X/Mtfmp2B16bujRVKT3DZr9UHWtSX/+wx9NXJUTLFlviEvV
myTC19e8W98LoLVIzjhfEn64zmb1vLbeHMFq7IFxp81hAJgn4w5gQmCIrmgauZJ3FXZ3/qqfsBRO
4S2FmAEqVdw0neRvdr4Clwo85KBzHNBHp2Jpzy8dviSZmvR9w0RNMEH7inS+He4NKyfzrAWgfDKb
4MHVFb6pslXdBOS3K6dzB8PdUJzJLYWueC3JW5isTpWCStm8O3nJrGQdoW5zRwjn1yXWoGSytA6u
NP8Y7yFh0eC99bvrcUIvxCjuCsd4TKeY9DiCjwWbE117vBqompcn2T24UkWcl8Kql2yfrm/5S5Gc
gqptwHkJVktLWniSj+cODU7DzPYHWHlhqyWrRWCl5ZPGRP0XokhitdubkpHpnK8icQG5Qhj/XL6N
hMyPqePsVtI1FA0gqA7Bt5Buv/rXdC/RZq+KeuS07SrPc1Svp8WC7dxjCce8l3alVGp2ySPLqdb0
1ZvV4mfqSCbJwOulMWPPQ/1HL2rJBWAH9Gtlj0MsbgHAqh4F3z9A3Cclfo4QvcrEIy1CvHdt5ZQM
drPNTHvwAm6Qjk5YRixR1cBMhQIxUmfN+YVrTPoH5JS0//WXAipXvorCWuV/dwm/7n0qW40tanCu
guwqAoa0rqUho2r8BdhOHM57IgTkUpHnavowENC0GYgrIOai4o4V3kFjF6kR92PVpuorM10sxlr2
NNyeJ2I+tCl9xWcldFh18At0SavzL252YzRzQPk3vY9RgSACcQmTokDH3tQm7vkfV8KS6+9Z4i0Z
No6FHjNIJUULZ0HUUYiuNElThbVLV8QxHF7k2aT+w/0ZjlLqkrioR4YJABO/jeEc5AkdzSFDGEIz
iVjINa7svBPSQUwJvskHoL9uGNGAJaKKtOGEqgY+0nKJAvBoBVFf4oHyvSjJOA1P0v5VUgfPZb1S
s9Gh+I0W36GIC6NNBv6G0fO6ZlqmaQx0YC6Hq83jarJ6lUTlyFwvIbQMVKHMWf6vdsU255MRzoCe
khjPChbBNz7fLmttcRZ4zqRlEgoeG2NRmZvTe7YHC8mbwueeUrX3IxMSlx2YjiApFwIdVGiLUz2o
Yv4VN1TlL4eW2qA26gGzhGYamxSZIPOr1Lcnn4qJHGJBuUgi3OLBPTFVjVpd9+8bNY4mfrf2nI9M
3styLV7mEF/A4BeDJoAQx/cfBXkTF/JFJj/n/lh6xlUW88lasiIwMIFkS09e1DaeXFdngkYYlNCZ
Ebyet7syh6k4mrKv8oZhVbnGfHxjL2h+lV2G7L04gOrNC/X0wXHBRj44UnlfiNc0yPnoiB3pHi3K
4VpbcZlV87pDK6ozZWSolNHQNKRjX94rhIzkTisjDrJ/ssDrpMNqWwuijgrIzIiRrqU0BSTAkdeO
3rCOyjtCBDvyMqp+VNSnholhhYGkGvFosV+RBmsIZMlkxYRpvsEsnFLOpRIsTC/Tp7dW/lxcQE7n
rBlt1an5FUljx+7jbBqR7PXDnvVayQpPTLrhtPI9LvgGf6dYswnVrHKpJPvYFdOI+AtpJ/uX6ihP
fG6nw6OceJ7Jkv0IGp98ccR/hzrn+VH6uiFuPMxYJq9o3Hee3cERvaubGzL6OE/DBQ2NNjC4vaNm
uFPg8qOYVI0LPF2+yFzmIkcUsPFWjuF6OpLmWeRg6gSbOcpr3QyC4s52+9p8uUyVWr/s9GGYs1yG
WL7C11JxXTAjWr1thf2GnozY8dTwj0Ut365NC2T5hGm/DE52uxqDNV9hbeFx7lghJHlKRmYAnhY7
2VldnKuLWgjGkhEUlIwJBWfUcPRmHmHgUoCJ96lq+UHdRNE2+F5ui8RZ7so9f2n5jINsqapuy3cq
v3BNXatB/miBVbGvns+W5qanltVRxTTapPf/qnNT87JVk9bnM5eXtwPWHuMYCvTTM6HQIDngblpE
iTuT2IUoBBSnoVKF3xALLQmtq8HuUV0RyBxcf5WQQbKoBXmaXry8MMF8Nbb65JiK6Gm0apF8yYpN
YRzezQUhej4N2059WgC28oGNIjBJ5Am3ds2wLpDhR10vFEV0izCC5PJZGITwBghcDp7F2AUX/1KT
LYvLhmnbvBQ8jF7dXGbxfKRf7ir5U0eYH+xaxXt/m4Mv/ua0VpzEXiVTVYLIRUUg3svpWzQ1UPMJ
FwMAB0ExXJbl4GMEa6T6mhOIEjIMt+hB01hDBym3AjlikElIV++7OOZMLUgl+a76QmM/6tmaMz2A
qtHPEmiuBNYc4CiIRgyZGC/hA1uNjfpvgB7BMMRi9jeWXowPSwmD4xiHkYP6olmSgVHmIMEoCNs0
aPVwSRgvqubhjbTC4GDTGI3c4rDo1WPP+rq1ITk480fDT06dNBFC6SvoKh7RL57lb/4hcWc6aTjq
N1AkYVOUzU0jKnio6qWF9HnFZUHstNHlDLJ2eX4T1gCsAVh7FE184Wh3tvvy9FHwZ57J8DsR+F/c
3Lu6AzCi2snnwqyjO5enKFaPuSxI6TSzR8X6mDBMdVYLqF9UnQweRLiWFwV8q6vCyA46qU3+edbn
pEiBWHnHfNA89tx05RfSQQBA4+7p5/EpuJi1foFHXVjDigQxpLJCnvltGCOFe0ZwtVpLEzMXlK3Y
W/vIJD8vPW6kAp6GEUAZm8Gbu8EnLHZZAtRzaPJJGXzutjgoSedWEOQbuhbDWlN3fAD4w9/2414/
M6KPKdgAuPhsPZiUxBw4PUPmPdxIT7xeKD3aHJHtG0ti0WhJvCxoPDRtfk4m1/CoULS096Lg8eJm
lvrFQUs1kltSxfvdnKcXbdQNzfiWurMz13RqTLHlomDif0NzcF7DNCxmZCetyQ8iaB9oUA6AxPWv
hkSj7vmM+bcCiMOvqf1NH0ivksdnWMD2nnEJOXFVdSfZMD4UMJnJX4Zfqlki1ZAIdwTSSfhCiQTB
+w75OcDbcmgSzJYD8UgFsDFIzoShTy/lbstXAVEF9GacwaRdwMEwzLXm5VsQ443PGMbX2l8Bvkfe
6Tuksn8K1prBTWVmhCRcjL7+SIHWHegIWfJO7UQlInef7MmvwMsZ11vy9ddDbgUQFNYjtXMF3V95
P9dq3g7hv6AG66G07cdTuinQxYx+y+JEPtwccGCxUo8WT+F8cD0M6tPHj3njvQwaPa5K+DwAXAby
GHBmDajCHL0UyeRTbSfI1kNqY6ZkgURkx2HVZ348ivlWWJAoSDE7snbLzvJPHEsa8R71HdFgzuJO
FqwV7Y5iIFKd8eIHSU479I9kr/A9s5GqOezQ7SCUfZGBsdM3PMUd2ETK5AVOxpRdwJEXb7WbggbU
dFqEfK4s8b5mm3h2ffc3rL0fm+IF9EZA5tXzpTaw/8J2OcYUDQGP26W7WuTgiiLAnvxm+BZ5GsqB
58oHcY1N0tdeqHmckPs25qdOZmXlbDBJkQg8eba6RTGxlTqX1toJqdjLskpDiGEsPzPdnzclZtt5
bKt0fhblwl1IihAN8Hbb+v2WFNK9PMlkiTrtO6mfdCo3Uj54Xd2qPKFq6VPIyYttD2CkE/fL6g3i
w7DJWNb3cnd46MgjaIoOfp3AICmKAc6HG6pZ1eIvRmvoPqOUJm6Hdkr7Cn+C99Rou4cc5wkLtb3+
GY9YIV0/V0urVmDzmM5qDSKQ9wGQL45VFISTIQSOXjkzmw8kAlgAsF+xIj5seNL7wZFvpLU+92Kd
BitPDgsndmsZFlMUwVdMJPQQ6zyCtjWw93FCXokz60IiFKf+qyaQ3r6JiAtu4n/BqeotuVAn69jS
eehKkR+gteAlJbRmDErBumAmZf0FqT6RDKCJukpEwvUs6p1EkQIFYXJI/YvWDVHaqxKFSFesNYIB
CJZ5vMwoE0WFbNkZFqAInDTidx+kEcVIAZ7PKvNgyW7WIvgvBlcp5q/RCfwBqndkIsr9/5NKDtlt
pZMAQtNc6ReIF7ubdWwqp2WwYhaZ8effawBpvsEiufPOOvQQu2CzX3s2A1eQeV+orY6ey+qCu/NC
kS/6ivsZLEE7HbbdeYtvYBDmvBmioKBQPEGiOlO1jjzsVdGhtfnnQtK2wmKPcIVKaBWbat4l9en1
v9qiAJKGA6eE6eWzD+Z+KfCTNpU+RukGaLtyoCyca8UbB9yssw/1yYl82FhSvQKlsrKXInxTwcOv
HbGErkX7u3yDKOroIpGvPsx5O2bK1QXBxKolqNT2Le2PulkcAHUIbuKpFV6LERfBQCq9g3uM+bIM
kCx6AWGEG1BMMO0yZgDbbIyCi8nhUJYBhdH6f+5i/7XZ7STNDeYBhN1SyfvPpRboxwSLG08Mfr9y
ldlTIBcbbNFQoeygcwPJwm2DGWXRUD5cHnWLFA4yzfkNUo85ka8dTGpRv95LnwHzWVhkKnn7n3TC
Z3SAWEXsnfyqJmn4jw8v4d/4GS5A0n+dwkFHGbQjncf9wL6sJyCVJtIohUgzkzKE+u7aFWZCUa8p
awXK5GReH4rP1wFZJwgKUd8D2c6f4vPdJLlvD3rpxMVys45YAjZch+W+jbbVfrY1lFNI207NxV3k
2APymfWSuVlO0vB65bCiiq+ZQkkcx16jxhS6YonXPHx8ke+ieWz5XWeTdhINq6acfmjhTlz+4vJx
72jozZTUXZ8y2c+aQgS+hwFYkgJNuyrGEn9gYhbr7tBhNVcfrEdQp3luzzlw4+MrLb+tg9hMI8ob
7S5PX2CQRH+H6mLKHaDIwxiX43TRsajmmdzZy8+c3Q55+maVUTU5paMjh6eF9P8378Xywh1mxfGs
9aXSOKJtYjR2+ggmcvEUSuRvJN11M3UHB3KXXgn0+M0fcIn7OkkCOzpOKNbiWRLzkS7uqOqveNHD
DRZImKCLAOlvDGnuJ3OVVcuhD8tzeH5UU71StKO63qPGzvX1RCisCb/R48PShSCjSaE0c/tLJmHy
gPzb/WahsI9R3aEVQnWx/p2gs6de3F0mKaiqrPLI7wAifGB7V2ijjFylGqGweh/uTPh9rxnYoRQh
HHPx1EQHQhDo2ArBD3ia7WqRE+0Ab5WUYnA+fS/H0qv5PUiWGZQcHaBXIN4Ld+Wgu53OqQk8GSLL
1WkD8cwww/iIkuvixecIW0C6KLhj4hgxbZufeF5iEmCnCiim1SaLhNNh1d+fStpWac76YyMRugAd
LNQ/mNuR3+U3Kp42lzkfTx2E+CZao05oITWiQExbHNipjdx+JWQS/UIdyWh4tO8qLfYbaC9l8VoT
RHrrCPpr9Q+C2Tl7lUT4OOmP2gDL1b/ss7/9vkwHc/+XnC6cNeDgkCyrOpSyioDmPbwYFRr0X62U
byxrLdHmMaBD0KOpLe0k1RaQ3zKV9DybPmcaUUUh0lWtg4OgpRJ7jAVhA9kZL5NpOwUu+eE2banA
KoNa9XgDGqDq+8wUPUiVjA6tNeLRcKwyQwYZzLdHlVEcthjkBdrcTL8bsDE4fQyoo/cchYarau0m
PTX8QWZCdz2Vl1ZmNkATHv5JsNaO9JA6p6PrVnfy0S7XzKLijfouzbJ42H+CbTthXgegJptTiGPb
uG1n7mUoz2Yz7gbAjrbWfKxGE2HtHGuuD+HuCJ7rPB/z2lLLCxe4P14HRcTarjOQoSozn/FDd4Ji
agSn+fjIWIcxghmO19uQAcHswopjg/kLnJubjWjAewIiHrRETQ7H1KTQIUj5DizWesW1A4YCohfA
FLsEjSDcTn/FgLZrAV3hgAcS4OW/4tVusOMtgjZ9XP0rDuL36Hs71vutQZteKQGj6dhhiJq2LEcW
/i4ce5BaOyzOxSUIU0/ACzlO7XKzsWTbNzkMJEE29aReF1hquIR8xixUCK2PC1EaJabEUI7PTC3O
8tRSXOQt5gbOj0TiVE4prgKAnfo6I9HWCJ9AtFH3T+n9TkCwzs/G/ZZWUn0z0oWUumMM6cX8u8rw
+mep3seR/DeMp6I0HNffFARkZBZ72y3xGyTcgE2v1I+8t7mbHVgGLCs6pRgqDG8EQZ09DlmkKfVN
xqgYPUaM8nX0BGfLbMarJnbkoNIjgQNlbgveuswV7RI7Fv3xbeu7Yetzg4eTKaliKdDzgs4AhU8w
sTdHQCQrGfns0vW8OUW2Wl+gO8Id8L4xR4WMyciDeG8XSm6TPa6NmWaZqgLNvCy98zlwFytbs3BI
ou6ZbSGHH26c9YfFmvBZ6OrhxlHDOGpU8F+Q7jYD+a3huvy1n3DSp3jd/FpsGtZMoaJfg5+a+BxP
oiGCO8YNH9cGEQD+uI4TOb/TrqTxdoFYxUQSFKnyUf/g8l+HR6lBI87XifZWhDjwSqiJM9mdAwIF
u8vy2QjkvdkZvd6oiXn9tRc7teNaF/16oB64H6z61CbK6Bond6ineVIepfCHMN4ANhnF+62xLV77
J+YALcxPcNnUtOjuGHi20eES+eWp6laVmJZjY94NmSy09Ajjeu8eMabmLYI8/1R0kLXurRDlDZSL
3knJPJ1bINDlXK+Jwc7U5FmVDiHQNzOHyzDl9PCisFpjNDj3T6AHg97nNRk0R2TvvN5KThSZBXgc
KOcpCviQHj4Po0B7sUMqxxFh+RwVsbJRsnOXfbe81MAjI5p0U34GJBqyf0rXoX0FswOzqhN4Rmsn
RxQRy4G4qWxR7RaJQuaq8WffPC62OaD+DN/GtHIidaI9uw+Bjz89dx3Y+/kCjT3pKOUqHJSjXcYs
TioDHOWTU+U923iWAhLgogLvHPnXxDYqusv0tdgHmw0QTMZfVxg1UEGpGXcg1hs40jdXtzwuxVXC
FTZkdtm1VSbO2TSjD1yDqkBAJMg62j/6y9ZNa4MbgPuiPwOnNMmXzCt2swoRP71tUzOtzTHys2Dj
MsLMFVkRG60qr0Ojzon+4vlui82MQgaJxna1Ou9tTtPPluyXIGERR/PXb8+P7L6tgNV+9SMbC9O5
ivsPvpmQojnklhwU9t+3cw7/6eL7lUeHZzpufXWTiY/c3GyIvm+T4BFuvp7frNSHuHd1nkNbozed
Ec6shjqAaKtp4PLy/Cw/FXTUWzP/I9d8b9TKHb+ebP7wNO0JeBaXmWsIbI/Yc9x10fsbdUFBnVvi
1OQ4lIP2WzGFoqGDmccZNoP0x8ohfZeNLHF1svcP2HivJzwMtfeuNOhv1tWDu0bF5+X8W2lbXCXn
7gjKvRdmGnhEJcakUey9J3mNIbv2OurkXFQSunMD5VlfVzJ4mJrR+nShRuWsOg4/MFBx//v/qoEB
RhtxPlqdK1Vb6sOY6UsTcjeJHOSL77fumBIBpG0eR2pelJwv1hibKviyCUs+VbUKdA1gt84UPtvl
1n3Z95+6WI5IOMpb0m/vu8+bLIq41ufiIT2MfJLFj/Z0FPDDgPRPn1qYHdDeFfW2YSU1UNBkAeVI
H0yNTymqsmTCsi6BARcvXg4UhOwQqM/albx2arnfR1O5Xw+MSeoJRCByMlBT0QVcgWll+2ny5eST
euW7MVnpi5LGtXiSuVcHSZMbCVWGe5CHNAFJyhqQyTl4BNuvO5XXfdHbVbRoGYG0sZAEl/8ygL60
oqhndr332sdsDK5wsVuvLRNtY4ojrp+SRWQa0UjmmDbhiq3OVq5lrvTZCE3ow0F5OII3p20YjiHe
Jdy2ug2HZIM1Oysyaidz7es+27uhTzC7Rrg6eBmqqbJ5aAfvfKZC6E5r4ao50hSLXviSuvjrWAX5
ll2BQxl3HTRtgkOoUXgVUQ7N5PReXKh0pv5spEv9DMhOloGsf2qohCyCdaXCjXVCzP/GFeDxRf1g
wDZ/msmQruUpRWHnxiVvN/Shjbp9K16EQSxzxatofEzkRalcGj/Knq6mZ+uFjzXrXY1x37uIlZWQ
dkJL9DQXvk12AHHe5ZAizQgvrMyacFGJmAnlBmi4/txhM0yXTg4fl7zxF+n+D3Psn+UPXP6Ydk43
GaISXoCPatRdR+WaGigcEDTy28YHGdUC/9E1EesCEmYfQ3JqA2K9ehWC0ecjzcD80T+rr79XWvvi
KzVFxAfByBDhqRseyoMVntOXllbXOATBwfzYjjvZw9n0j7cOyNrnOCyVy/PSL8MxNqiFFw7P7/T5
3QfkIy8lvSPUW44zwdyLa9mLxZFxPLfhr7/riaSYeUcFhq4BZbF30C7CNKn/8znleQMlB9DE4sfp
Idgajzjc9T5kHLZ/wBH5YJGDKj61EkxH8sDhCAoHkW6UEMoZM2QYCiyIpAFpKyeK8W1vrAuKAfOf
8Q11/ybYLvrXVsc1WVi74cKjcM72HE6bE3JSp1eBZIU7FZoGCbBKgd+RXbHg5uIhubAP9+EO0syH
lxQVpxwldhKCRk/qfhHeP0+BiY5fmISFdZ6T2idFfJBhwbcxBqX60z1fK1EZ/WNS09kHb/Jocmfa
y40ZmcFZvHn+Zg7KGYb5NOwWAUjoE/joPy73MWZIMSazksQDjOkH82WH2r2qiWyptUTCe5fKHoCa
PA3u8CPU0uZ2t+BOp8W/Ov+UZ0B4ARc1E6rXGwTevO/jwzMhOib7+kV4nDWbQkYyqE8RG236cTmo
+pa0itSl9hPsbfWs23ArhYjjgUO66gGuIx/wJuhExr+G5hOvJnuPs9OrvN9TNQ33zhdLmiIOyddL
7LIOorpC0u2vfXLZot6rQEYGT8FrksYBnT4IGHWtlUxY2rm4ETExYCo3OE37tn1TifT6pVasVZnI
2zQbjv4+eT3Z7IyHZNmtubvzAmCOx+Q2x6UthtZEhj5IyjD3JlhMXs5MpukpFRqSqOZpSCzvF7ge
OTYaqLpvgDbkJAwpVG4x8y2wqpYfx9ibyXW+maXdU1x9HUvLRdHuGmrK+fmw2pKMbptQqSLRW7BF
bnwywqbXDBdyk3SQPZ1cu9JxarAo4NWml/pGhuHI+M0Y4TQb4niA7RYVBzLj7R5BFgKQwFx135m1
851LsWk352BxtWs504Z/t5RK1820C+dVWZTDuUppTkTpZbPfBJsGgVFNGVoCa12R38YOuC7KeZKv
k//myZVcQRmo82EFJwAV79MKQ8MI9pvYZA10c8i28xnTLyNA6aS9E75Y+gpa3qH1nTwFHuKlez7l
WlezWPShrLpTYzPguUhMA41wxDKAxjXcLdVjFFP7BFmaQtiDgX4tHmeSdlDRG4eH5Fp1yi0qak20
P0uvLeJq+Q5nMqbUiqZ0QOAZ8wltOoqfD6lPSNJ1YMVJ/3MDaJQ1y8ATyKU6UK4qjmjFSr7JEia6
81n3xAp21sVzKuEfoWrnJIvB0fVjIFckQRTbqEwRgAWMPQpWsN0bCzYEYjMv9lDwDckpm+aCKe87
egYoX0dBICL5/6eXn7Zc0Agom4wboc4FAdgGNgjWXkh9Ai1KInAyzYfQt2HAKzuTUZR96Wl2uMyW
X/jm5CF402RMpX3p1/3DIFbcHT5auiIU1YcyohR14DrnLg4AqhPsnbODJ4rLav+fvRL+8jUm4WWV
+ild8RSnWEnO0RFXfI8JIsrg/FT6NrKg5DzTd9wgNk2LXmbB87FOTqcJqgB6fwfRd45w8Zl3S2XX
QWJVpgg9+FJcW/03MEdRrVSIHckBxmiSrNQFpTJ7S441sc8pjZiJc3c+SScknpEUetkLFW/1oYVp
vAhQcolpT6sjWh1DJKuPpp9MUxLtgAfnDDreALpw3s0m6+x3uOZWfgOQ1hHpdEEwoc0TODYG/xSo
2g69VNBBZTDGDWYURKlFs8Dy/9tZw6zUvLV7mhB+mgO/D4iOaoLAP4f04V87yuQgipsaky8C4Go9
SuqJJeymd/VGlhVW5t8I2NrVeDBNjJlYjwMpm0NkIrKoLsH7GXGIz5y+qgfIU/TwqVoHNvET9wQN
m9ZmaUeK7KSe2LDE0dDYO3SAaZpmOfCYctTrC3HuV/bZXChQUQm6uNxJn9EpsWKSskMXk4Kh0AvT
pciapzoWSaAm2DS8nyTl+SyzloAPnglM1VkK+LzRUujtBmj8k9tihBZJb2NknNmM51Iyk3evR05M
ejW2daipEphj2CLH72BAe55Ekq3Nin0EAOI8Pyho7pY1QlvCvtcU5+92vDnVwhaiXtRhEskAf6uH
r6UjtibSzBkrTHqCIqev0DQunUMaE0ugd+D2Jb9s8XvlwMBo0gJWInEZkSVwv6pqTWHmsVTDEWer
rsdalTsImKgExK2ucpPUX/gAnYN6osUklu261/vUNDkOGRMAZQMdMx7qwe7TnWXYe6CZX9m51eyk
wQnisLOSi5zHocnTPDpE/355UhVy4ZZVtqNLI7gs5FEOMnRkU7xSVNDYUwj5HvkPF2NREtlQyafX
V5fFhi8hcNKt5PPyZbnaFZ7qKqtSqMhrhPBsuygcQU5J7ROAvkmZOnJHkz20JTKBbqUISHIzhiMx
hvV88CO5UWIDZxLwB1ZnvgouKjfAu8joDLGHykPOMMBqHcsnRWFLPOdAuv9G4tdZLA9ee+2xwtVJ
k01tYBbytll9kKI65VzJJs8fdX/R9vMEallXSjfaluw+QP70PDu+Q1hIpTzDfI7uQ8SQcGziS7xj
lL42XaJiIK6iDCFO8FLtPeB1ixuqLV3HTvRd7O3Rwkmlnz6NfqH2ywt13gtRMd9xhYxvJFe+pFpY
3AshlWQIpMH6x8czTzIII4sy4VLnrzm5eqUCj0MR6u8wqaRORCgmNBMsF1TbHsgONAzNP9MnVnEm
aXngxnPYPqw2+ykjWIxXSueqMxnbARbBG02H5Q8gzLf6RonIW2y+R6XaWlsNeesIxyr2b3AuaGXq
8q0ORyPn63Ya68mDxJa3Z4Ht0p3TcLfxHoDNmLHAuZUMjvTmSNPnP7xeGjJ7PX7SF13pT9IdVP/p
aUmiEmZs4mzt0mB38QJ/nOnTi1BvZDyUiLkwW88f66HTnSB7SDczeCAvWS9z1R5qb8m1IydKAVt4
AB/8QnhSjxLRC0zcAz80TrrR7SYfIuzypV7qXwNRAqu+A2ULnDzQe2sY/VCkYGyofgFhBpVB1fmA
3jWtqhudi2zCllamdGPkCYGBWSpRMMt10XF7ODkYcqAtXLOBsKsWffU2n3zlFilGl5VcH0+O+0wS
HsyxDfadhdBrPu1/8P8mTZlSoAg+pBv0H7lQxcNQMUrMRAeL8kb32kLoUBbrD9vuee+KxvW6TVfH
vQfXdQVhHQ0+gq8s3pokGf4e9lFzocB43ImRigZQ64ZgTpKZVuXaUETKvPQyZmFewQmvRw1UvabE
BVdIT29NnCBqXouRSnEKXrrLgNQ9hJfiEb688X4Gwo3jhr6i+b570olHHuo33MrCfwUdiRY05i7t
YaRaPoGkAp7TAomCCRcLpArMvX9s/QguuAkj6yApg0lwOgaKPb+i30zfZFucwSV32Vul4fa8lSR/
0Cy2qczaE4KHYE/7xZiIQVxTQ7HUA+1brdi0zKKl7/AXbjMA5YWJpkB5V+L7gZTPjYIQaLVMyt9v
4ZkwHgQ3HnIFbUZVKPzk15l47XG3+Z3UURfKA3D3/A/LY0i7Thfbjg9/UmsQrJPeYvaFrbekAvQC
6P+B8FK4Xny6H62yWjhYqinwTqQeVylJCtRqqmKhcRz+yYfgFMz5aLW5LcQmAQW5xyTjfwX2m8UI
XlowBMwb/jcuf/YNOA+wsRTAlgJ3U/Vpe65BYLM+JdXcbBi/e6mXPGPWYeFtnSgo0l8in6GHcrvb
WBivImzKenp5KK9bROrEHtwVxPRIgc4RXLhgMdydiljG5amnfN7ZrkpqvUIEgoR8NqYaF2JVoH0Y
SdKlfFtNVjixSgbwvSCMH62uWDgMftBypnZiTuwsCqV3pjHP3cySwo6b30S8/2iHPQW/DnrC9FKd
XfXJB9gQgHISZvdn5tMhMw2b8eGGd94DZ+kSSdS9Y7QWFtklW0UwaWw8s6Z7TUXBBn1pHMJxt2U8
0cpZ9m8cmR7pcbeU3kAA4rV6gbBf6qBQZHBXyfqMcGV72MZtzUqEECcQj5qu0w4fW3Sk9WMPclu+
DlwSQtOlR3UfeqipE1xqMEoQxbjzXJFBnMgQVBiUKaSGhHtJ0c7civAOtQmlOh/ScTwsh98cHfTz
XT6CEZ3o7qqncvCzPGj9t1TN9ux61aB3QFoZwotakp32dohLTj9082b0oWDO63HrN8Raps6VUaHN
AS5gxHzpzC9gcCORCpRE9Xqe8m8FSYFn6qsUJWhnFYl4wDGrAQjoiwrKQ7zO86JIyUUbNHvQtf4e
d5iIsHP/KxoU2fnzEq0TaO60mWKxQyu1OExVo7BsBDhzXwaVkzdG2rMxFlk1RhXRoU8amS6W20B/
kEAldQosOpnSwk0z2e6/oo0zge8vzAZVAtFPYWt3NnH+GKqrQSTLr7CgL/8WB1kGYufL1sT3wFl/
SqncH2Ev71BCQfB8cC0N/BY1ZlDXPIrXtlMruwIIHLYX6bbXdmE9wihTcPOOzSpiFuGe6raVfNWL
hj0Hi8BISqCr4L4cbzl5XxxsKZMAUfXVKQ2pOBe/zVkFTjhq9/1hyOQc5xcLYwMRwmTonM5c68/Y
RAiSrHPWdskfK19C95/0JsAmBHBjhOMxh0bhiX6U6vgdEzPMtkZItrZNphFP3ezasQKnWxtqW5Yn
5XY9d4d4pHTIV3fY/UhtnRJRQJbSfSMx8nlYjThRur0wn2968n7IZoP8Gsdm5306ZU0XLSJdTnDR
oJGvTkr9pSH3sTfRW+kWBYO3QxRiR1SI97RhXhomkYliEbB/A5EIpZkP967qUtyiCmOAqJcRIBdX
/evUS7QsdOakNXdJgFqpN10kmbWK7VAssTN/tiOCCkXvi1IWynZMGL0dGiz1h0apdl4lLgAlAS21
bWn5mwLfb4j16bXLdeSTEuaM8Kmx08X4gdAlmMEw8w9jXDoaUBfjoMbQ+JWWcedKE4DIGfAl+m6z
C/D9lbOsL+ySFROXnGLUyfQrUg5VGGVkM7me6zDRpFRUta/KYAaEvh6vp+ou/8+xpkfCcsb6i8Dj
RjodWUsXzcLqAXMAa6WVnOxEwoKB9Fd8eoNcHkaags9E7TircXRo/soVpeP5+MfS6LYUqdqbMBIG
B3G1mQ0FQxmGvKKmp4oTH7WIKqhNOeGAFMHsndCcUD/jAZaSsWlAhxdUJjbFk33fR4TUBqOFjI36
GwuRbrVzo+GrxsBN8gln4k2PWOEcCd/N7tLN6NBHoP40u0DltDSEYbsc7FfiDz8x9NIdlXfhtD//
La/KhEZhOPk9X6fCSbCWOHoLfBNIIuUh8Z/BCVKpKyBD2VXD4Dw0J09BQmjWo/qGZFS+mPUQlI5z
6/FIbJ6B1UMosAc+5HhdaTYqm7fRn1u0g20q0PlYnEx7zt2scBP3WiYwVgDFBJ4/uEZOOR6E64hB
rRjTzW5Ir2nzBvmLhjswv4EhNfTD3vmOd54En5Yn0xPen6dtyfeiq9USjhtS3MCsdK4M8v+E0U0v
rpoyJb018mjagjqgRWGW9bJrCXKYThrEmvXYc5/P+NfWc3lCRKSdjLCAKxRk4Iv9pXxDNwQ8SQ3/
LXIzuUhyHZzR1jArCeoOFPicxYpPFYWdkAZ96UpA5gR3bmXrbsoi3q3YmKCF31awvW87d/akzUrK
MfvtSzRoab7yQQ3V6plkKuXqjdK8iDuknFb3DiLqyl2AzCwN3MGw4/PDj+TYHYHWq0nhIahHZgLc
QWyFsuersjeKl217+5wQ//DHTaOWrim14aQpUL5eyNKU5g3dzgi3oKsuii112dG0ZryJ3gZ/W0Es
v0JFACCpHQLRy1Xf1uNnGjfr5587vZaJLDnDPK0bEK2GiTYXhc9mdXRAvhcO4aBDJ6DAwyObajoa
0Rd9EQa4p0rxKOV2PQdoFxhv1ThU1Gz6iDxMMdmn1mtocL7jlFVXZhba2IiD360dilRZZcoIDO7C
eoTTA0/HpHkA7t+iaTp3tC0+SN+50KZVlbTOXzSWPY/DI1hpAqrE9byDUbsX8sVJ5TbxsdXkdkBA
ObInDc2//hE8Nk0hL40Xd+5x85M7zHyk5JFEocWyHy1gd10nFtcUS+5uJJtu6Ldx9WjqyTYXjo/e
UUcOCQAsG7Yp/5BcB+OREvFVBPKI/kXhoVVij7vSy++La9pROYDCrvpdJehTDUMyv1wVCYK3n4fs
6rMXaOUTK+zcKxhB19ZXleuGx9rdE6nu7pb1PHUQf/dyrNflOo4XOj23HNQE3ri9Z7Jd+s2GLs0U
tJPCTOXD576h2HRhkY9/Pwwk8mFW3oVenqvB7JxJ/ptndq6lvL8y48pr0BSni8SSXX8bZV/QZMar
eoF3W7xzYlLEJgzgy6EgljV3Elc63GCuF3UAw8w5jeULwG2LK8QpJk5YKz6I4LYewfJ1X/hMsfK3
sW/9C6GelS4ej8Hawe2xu7JPrtB9U8WuOfT8nyO/C6sKq5UETtZe/afwtdG+Zw4nV4D2jV2yvFZ6
bgUx118hRV2O1FoAmwB1cZq2SKMn0aUa8BPSmJ9A/EanyqomC2KxWmVEyUdaGWBj283iOtHL0Ljc
AyX7LQrhfeIiaLH2HKhn0doG2Qg6YBoPv34Z0VQ/uVWUeHF0KArLCqJW/wFKfxiHcV8YhfIYyC9D
6+aPMdC9OAnZzk86pdyZeUnSFnm4Vx1p7MSvFo49bLbEA9LPjlelZ/qIg08bvkRlcmKyPHuFwq0W
PsTH9KrQcqKyzNOjbVZvdE27D1xh6G9Wwx76SFPL8E3jPoS53Yw7grxzCCWbUS6cDjvYsBMPgP8a
POj8kSGxyorDVZL9EurfDVa4sAId6PU1FuFDb3wFQuD43AoezSZqKInitx5ufZnNkOalNHVpQobu
U0li9LoSU97yj4+whIQYs+8POp2h16isflN9GERVctZ5JTqP9Xvv7C1/RUZVnzRFKvvgIsidEp3t
hHNNffUf7lWKMSvhvom7Jp3HIHMsokYJjFXCnDvFCkb8pezqkJ+ArnHEZTUO7qVwjQhuZD1fH8hd
p84WXLVGHNw+IFIVjdYI5giToIHAc49pgvvNGEHaGJ2Q9sXMpPAMqDA0nVOE3hWL9kfwRfh/xCcv
5GfE+w3xaNGqSM5iWI7ieD/qbvVeNRQ/4JRSbyYei4DIOPiTC4E1UNVPiiopznHDY6De3nd41Ggh
Uf11BCqbB4cIgu6q/wJCSDXWYZIrFE5VLRxvkU6l2F1u0BrSy01QMIshgl3DoUA011vn5Ks1T8hK
8t+zvuqJxkzI/mw2v1wYA9ZPk6TugHD04xPjsRzKLi4Rtm+SXxk6KP/rOfM6qPDjymSp/epDrljk
8WosWXQnlCyNw2cAoCQ4AXItIVO63MBSpEl1swSDrNu7vrL8kRepGH2v4YO41lk6fI4LZdwsS4nT
64Q0qelfsDw8Z7H6w8lwzIVwqfWf5bCNgJ42vLQ4P2/nYey3h540jTbil/1vfI+1zO97WMdUVma/
0vVd7LkWQEDB0qHKebp/5ybs5OL6BgCkmxpOgzLFqwr71SE4atlPGfUskd73VJowZ6d06GSkjLnU
PT1ODPguCxYVPRlEA7sM5eUPk4MJ7HVXRiG5xZ/WOTz70uFcFCLQo/eLv7JrJLbsIa//o1HkUnOD
Cxs5Jak2OD3UwcnYw/GXMG9WC49Fp4JHpw76kQd679KUIQc6J3RLhJBE9/GIzUw7f6JwZ42Bn+sH
5JiFAK31l0Bzy2dkcA9+hw3MBWtr7adFQR1iw6TNnrUDpjdBWToSYdKRkOM4rbcQsEcvUhR4BD7u
EOMxhrqxn8lVV1qf4zbTXHlXdF5Hzuf+mRvPmaiDWoiYuQNqSk02WGWf1AfCYGIKUnDCZVDF6IRf
J9Iu7lmX1065WkDPxsfSq/Z/X5Mz0QyWMZyzy4Refs8rs3+L2Tym3CMWEtwif/91ACr3pzr6AC/m
k7S2m+UGIh7FJmvuQnaTPYPDV1RvWN2UcbcUO1O+DdX72o9LkokvjPbvMhflxPc+nDpooAXUWhlT
lXV9Cgq7epBae1Gf2xuz+S0qgx3ySgh1tcg7FnRzNz+ylYuIdfGPpG7SGyDSnNSWvaxGZivn3e54
ZO3potaVZw1H/ENC10WZHZ7GRPXiY8KBE18r0Fo6laRuIfR2lyPVR9uOTIB9kOAvtZH24rx9K5B2
sO9sG35SpIEpVN+a4KHZZMVdzVu1XdbGmuf9Fwm8VxkLwSjthbzGgjmI77G2w5r/kyznMiSSY0JP
Hm/ZJW3O8OwrKnTUXGuZG7CROQW6qM6syG0v/6+TDPAUDm2AP8ZHEVd9+oCAPLft5kdKsz6Pz97b
zy2L4QTpSFOnJatQE81vd29A+lq78tChj9JfrN8g/BGLWprDPO3DbX0M1BzkJxVJpYW45LrRRPDX
cvmkZ4pe89Pz0qpKl/q8GHcH5QIbcOuEY3rfuTkljVwjIMO0pOKqQGKMWtQZbEIe7GEUjt8mtQmx
ULKfgT22zTuG8/NauzseMvAplrDVqzUY8zS6otgQc7W7CnNAjoBJ24+3G/IAZOVNTnLSp6qKKynx
qylfuCofcRHJ/cIREN2VJj2jIzAWuqxRqj+5QKQYecnui9PBcOu+tvF+P2QQPttjen4SVbenFR8J
UMRnfBksgAOMcoV778eSPyRD5oT5o6THCrOT2N4YJtSDMsvqBZU7MwfuOQPW9EaO+6E9mrK3p5O6
BXNCg3UZ1hVD0p4N3hUy0IgkPWXQoHKGEsidRCa7gi/FQR6NDZ/y27POtVCmbDo3+gQRwnKBTmBL
YdJbtorvIkaiIXJkqxjEXWf/yGlpb8Lh9v+QUSYTE+GhZvUF21mEAE/XX3inQkSFf09OzU18CZ8C
BisN8qWpKSTJ589g98zA5fQEf3LyzINWkgrVQZN7+V7gyR3sFihhpGcrdmWL4kEzNImRSkRl+rTE
Pgf4AhzGhRYPicQ7hvY7PYA5PqnSfIJmhpCNiCmSSFfjz3Ns7STsG8wkpRMCoxzKPWeG1JSdFjbh
wEUQAJtzDO0VBaEZQSngBUC0ixuhTMmSK/O85WSqCaks0DY/m4ZrJyYZdo7fHRoP1dp46O/UDZPh
xqzL3kX7BsMLhGrpWDvFq74R1SNiI4EkcEBXPDKJ5ntpwxIpGCW3jQVFF3gOiCNyKZm7LFvpArlM
KXv/sX50xkbB47ltzBsKmQbsdVYOYFh0fn+6+Ht2IPtCNL/l83HSlF43IB6ZdZtHEkcI9nmkFqUG
+pCguB/mCM5S0qJhK4tYSqX04A1zmnbSTRS5T5BoJD/Sd/TTagWCdVZ3q1YwvKgTurgEbTZrNhon
YcKwBTCWi9NctdGEUY/ikvmhq3O2clqNEkOglnUvhQYQ8P3WOHpGL9Ts1hCzHwMu/h605Rq6bCWU
lo43OVH3JxkMg5jQHlgnZ4UcAYoDKEesXfCqzmU3qWV+HaworQ995uk7hZZNTzYCDYhfQ1fj4Dsm
2DRWKdtpJZtcNCmZDFktt98GbEpMz9b97xcn3YIF0GtQAciG1v3gwxQxFW0ClA9B1Jm0DgPfsj07
d+3u1WTxOli1By9tc4CNQ0+3eUTauLbT2JuLFEZ1c4MMKqr2tOQjImuwV1S8NgXjEy07p4VbFXx8
b2ZoT931PwWGGr2vNe80Yn2/bZ3uxkmd9VHT9E7GBI+4lngoJyCNk2Q/QgZuubeohIw1LbS/E8E7
bG45ZzxqmGShwfNkypMd7glST506kBMdm53g31iwQ5qn1FU4fQySEaq0NwuABw1feXGzLuCB5/0k
poY9DBNz16wYo9Qdu8UewrciOxZ3RqQgZskdzK+WflnTJyn8hlAQSzIzhlhs5/aIonzQFA0e209b
vStOCHqHVOY3yHNIXyA6LmsdtcjflKukXbpR7cRoTRfUdOnqgY7QMXl46ZNRo5N6mv/GhnREI/0A
Bzq/109XnQo0ZL5JT6MlHOm/Z6pTXhnLiiYskIxkTZcOtAu2WOW6EH6wciAv4vrvlv2cKUZEN5n9
LrsA3C9aVMmiO7PhlL5hWTv8Hz1EUCobVsbrcZIENHzfioUFFcN4TzFM50m4VoPU4XuG4+swN5dV
kvVoZABP9UhlF8+tNo25Q2Dwu7pWD8bHKRR0WzYr/oBVE76kjb+pY55zfZnqAQ9KLg5hcqZDNbNy
fKmYMmfSaAGzQLrxz6058z6BbyFHbFsqiLQh26wlkf2qYRBOa5ehHkA1CcjQDQlVywOgQo5SWLoX
dWUudg6qFvZnpM5GP+zcQQqdcykXcG1y9WN8xtjub9XPmyJoNfKSynSLA0zVw7Hr4SJgdO18w9iL
WXZdvjxi5AVYWAajYMiuSAqWiB4xfAJIdVIBBDnXH8TMXrU4pQHgAYII7c8nXApytzd8JepxKa/i
AnBbsIOa2Xv/dXiTTAqAdnMhk/rfPmZcsgtLHppdT2+mDNugQF7427ljBziUUde+uPIUD6IJ/d8K
jKWcB/UlsgvBt/ouJhYWhjr+R2AOCipRItHWt/IPDbdFGb8q8bCMUlDNA8/9HACmF8Y7P6t1pkP5
uyHy5RQSCYvColEyRa3iAPH6I3wBVhUY8IhDpNQ1RX/gN/dbLdvJtz717SVDBnimu8/BgfIpTPV7
hpmJTKenDe3saIkLQuXkCjM2+XYqH2sdU9Vq0JYnKuDsvhlg/pK5PysbeHfs6Uynsf+Bc/LCfIrg
hRp2ZG2/tA+W9yH3kiIGYLc6PTYLkWMWnEIwT47t96VD6XWp8y0OzQuPu/bABTXdNe1WVHEX6zkv
n5H8oIqIxVNkJSAOnE2u19AOgksWWPxzDS041mwqDakjrK4OYN1ySmR+E6XmcyPZwEyQGzloeA9E
N3miPZ5zQfbEK7A9g7gchgxITyhCJWUDDRTe9FKYYpwI9ZAVaqEOvcY82DgTLytQ+DQAcKrdSHEn
4/Tn5g5673sHes3q/wEHBX6mI5vZZEMyLCEB8PVC0Df6Jp1kLlAsn7MYdzxrbyVjcEdI/khKyxC6
yn3dk8m/ywWiOenw7CyQ1g6Bcu0AQqghpn3dS2IbFkwJKUOJSs5z9uQuLw463gQMhz8vu289IIW/
idMmYBbnFg5KH88zFaiPHUnIsMlrjk5O416W7D1IaIdiRU1MePDOfUlYOzaL/SB38j1Meh8+w5n0
AcLGPliuTaxR5qHMC+UsbIWlDBrpHO99+IJMagaPWXh9sJkWd8sC5FknBxgrxzO22Wz0r4ju3o6K
at4n8A1yKjv+YEYQ641BuP69n6kw8ba8qp7w/EtSqQOmfHLm+JVk5YIphPnTQyzqSCj9LniM3bgt
BQC+WxmfwlwnMgXapU5fIe0TEpB6s3ICARog16D2uwRdaLNDqFeZadeg04mvNI0Iz4FOpK4Hj5sF
0SF6EoN/1Nsclj+MVeK1yv1s5cY1Rm2CK/XAHSt3J+9NVplcjk5xuIhFC+V3YlDyN4NTvGRrCzOO
BUfWKsRI5HBZ5aebEHQFmLJpYFy39szY+jcVWyltZbjbLhkLfnMRtbQRnwy5z7a92WoT3Bv1lV6p
Ww+TPjiMF0VXazEKXjcC/+LLbRp2BDCixwPFtbDXmwbDdVRknxIk94Um1tIgsYkmbQpPgh3FFxFj
JkaQpVCcwuv1/BPXkJ7MtbaJ7ymk//GwqzVC+S8PNpgB9cfFlN5PXX2luqEmZEfJ49oJefJuOddQ
Nvs8Qu6iXRqo6oTw0Mloe5tk1+gx3dXK5XYvWUP6rYHRKcAhHth+Ao4Z/wqEJTRM9HPGUnc2lUZd
DNfUtxJurF3ITQFTh8zAVip1/fEoBHZbQz2Na/whxu/yzWEiaCnYFnu+tKAyO/P7gzmDqT5unkXJ
SexJJvqcny8prGWLFS8AZR/z6JLWweAxjuf7B+SW1MBu330kb1AHT8pVE5pT/Z2vCRfy1ZKyAjgC
xCdnZbI1xoEGZlfcMCKmaW9wDsuSsvPEMjEBX5pzaK7GFAnafBF6HJfL+SK5Vfm+9WTjy4MZfEKX
STFnPkxhWUGN3gPTBQvKg0lm52qK5N/dODQn5UYXsVH2COHFsbsJlgh0PCQlxoW6W/nLoGNeVOFZ
E7Us9+uGsFSG0u+e/MOfj3yMGHU6WBsQRbfy8ht+8HPRSTruDxkPNQEM3YRP/GaV59SvrqWLg1vN
HCvrelwjkwXx4qDrcDwZ6Q//BJOLrk7+0XWYbitSxB5TJBlGfLBjWedzI7TaRH60t+6Hc7BFFPFL
eiL4O4XnAypwmrs9tPwmDJaBZ1r/C1POMcFRPYja3aFQsm02/L7qcHaWl6mtJJGIvm7dW6hCd0vw
ezxcnVkCsctL9WsjUfvo+1GdEych+8VzTpZJGTf4cA5vke9l07q2JfJsheBMC1G5Dvk381u7MbSI
KL8hk3VSbmmNu5+A8JvNYVyhkLW51YCptbd68FjMY6l7P0TTWRpQCt4fJc9pRaawNUHGRt9j0WUJ
GI93k5JCodQZ2nIx8jdRf2Sl4+Vb0XIejmJYZ3PTv6Mn3skqo20fdHphlN4X4qhp5ZH+W5X/Y7J+
2YGgH0nZ4BIDtZ7esFEIoQgMC06/CaFmKKpQoY3k5L3vhxKR68EVWW7OYAcKNNry3kn+S+/rdPk4
N2E0ng1opzGqlfPQhb36oDUFq7lyFbaHF6bf50mqopsAPZZX6NQRmTlyp27iTZS+z9qQF0r5sGzi
TMYI6Ut1f2my/0G9ym2Zglr0PtmyZBv1KIDsbgDAxVXz6ousl/ud5Ahy6rVsXvu0j02ioBv0lgdt
n2Lm++q08j7/dqDQWfqhWvLGMt5Hvo7dCA6XAlul/u0z1k6DBlG2qPjHzcuQqvwIzT+GDsSBXfUY
JXH0DLamQtcphxgvsj0l5mTKq4W43XHzGTN1X7K8YfxIu8GwXNbjlTP9HmAU5802IfaW8ZnlRknr
5RkbaDqfVdQXJIbT2hN1vttaSvAudWpFt8gWnA4K760VJzehIe8gWMMDD7cRDCo2bbHeVG4Jajsg
eZrPk+33UJ3kgUGIDVx/0FHGNeqBaETfk4YZbQ/CBqphoNo4RB97vmQPrLCqJmTihyWwiq98be1C
qPFtrZLmy3uoO9xR7QNxgPmTs/FDjaxkgI9GAuBH6yXB/hS4Uj+spitLTEt03xfQOMFEGR1YxloB
FVwl33uCkoetik01VE9Z5Z/LLRokrV1zxxK9AsL+uScXEqu9Nx9KuKn5BgTy0j2rgi/pQVJox9/4
ADTpKbg6KZhwdwN0MZc2exsnj1YIEiZcZ08W97N8CdfL9SosuOyiMa6i2qEOAVMkBJHcIKSCg9vD
2zmCbTrGMf1Z9Y0aTEzr6xThoixUamZJkAjlb/No8NcHrkz3DLPAfMrcnaQfkJdyCpVd+q3N5r8l
44Mgr4wNXETkn4t6kmuafJx/NbLcoGdwc9ai9ZuOeTpJH2M4eBlfvdkaLz755aSpENBKMWj1Z8P/
LuAtk9e5v9VJybwFsDwcw5J16If8vrgKJLU0+W81bgD+H2IuMJQdXTeVh7kY+aVbfeUH6Rb/XiQe
CI2PlKTJ0YLb36JQdNa83z4FBQ0sKbdS9eZgT+lqEykTAa1pNRM5XNkiJlka8ElA0ytVh91tjg4b
7LIcV5OGcpA+zNa55IY8oCDxnWt+GDN8voj2CL704OToXRZXJd0vNLgXqV30unySj9y59IzE+tZn
1gtiylonFcwYjzZaAkXsf1X7PkCuKUH5rh09hP0vsXdR4DanFYf22SGvUYHwyBY8Wt2cdHTREJSV
QUN6WmRsxL5LAc9rvDvKJ6Pru5SzMyhVCwCCv5FGicvwXSpZUVk8NilWjV3jcZe3rZ3uvMYdSSUN
DkW+fREuibuQ2z8Pb2NDVUKcN1xNH6MAb7uSj+/V6xgpWg8n/nkqIiiZ0UCTdf7NUyHSSriUTSzD
YMaNTeibWvCrlqS34ul7NEBx30Qd2ppxrKfmKTsJ/tebHH+Pm5NsB4thDV1lY+aAERIhn2l2fO9+
TliUi9MEGfouTzXPxOLiYm1VmS84Ex3JD5INL4lqJzQInGcQ315xQkQXrPTXf2Vuhn8EOTRvhxW8
mjrhciHbpaBIQSzViBcoL+fnJ5YLu6quamR1aru5kF2exE2Wa8xWw66EVn+htE1QmQ94VVriuuGO
0liTq/PCXcD+Lsg2PFJLvYBz3QHb8R/gCMwk0i6rIHTnXxyJBFMddMc6szPGS7WLa7MyXSz3Gg3D
JN+gjNiNhqwDtSRZkHoJ/AB01yvSELRyAHe+EFeWswRY9ONgEHtP0AREjUMb/GkGb9RjQOgaFzNQ
9OjnAruq/xGsKWZG8XfWlrX4RITCEJqMd/AG2xcosIeJMaBrv+IwRznLt8X/yczbeUrM/fhEZ9VD
T+CQn41Rx3bNISnDOVnkePVpJR3tg2m8i07BHp805HiLwaP08eCtbzoAQ73Ue4e0BwoKBOUQgKFp
Y2goR+dMN9T1W6unMKLTjoBt7YDi7BRORipFa1A5TwvGudWCT2wWo6xlKrhKoLOm97cfw+Fkty+4
0J6JelGIMoSGNX6oZTDOp9AE5ncBozTeuwuNWLK7rgDdTQN86vXqBXfvM8efQuUjcRhhLkPyeucq
wPFNBI0LBoVJTgE2Jc9uxp6E8ZpROJ6ocWwkrL8SI9emykHKQuduwvQDbnXSveD5+vpqg11heitu
/BTCRUB5DBQUh90SC7MQwkGf0p4De5khqaw1nk4ircSMXgenRgmdXRueF+sBL/63AlCEwZXfknmz
aRDqT1WWD+Ak4AkwM1BrV+8fl9QGYPm+AvsXnivOj7Mmv/WKcchlP31IuJYX+cvTgzS6tEVPfqbX
80NGKyMk54cdXbR46Wn8wWvDw6BHQcWSoHwzn/f+ax1LNxNVUILlPQxVZvgVjoutSZT3DNoy+buL
FA5v31de4aUiyU5/Z3vl2eusiSafnDuAJ32nl18GReHsTyV70nmYXJ6tqRavvRkmoE9wf5ePhG3U
RCPZEXAT8un57W87AiS4LN/6KFDoEPjLfLdMPGl7u3+hf+xwIx6LpMlY/kz0AMeS5dWdBwjhXvMb
e7VLRWD55ZTF8FkuQBnVeRK8Zwx7gZ5e7AWYWp6OvX0SCRC9WAVxEJarI7/uZC2egbn5mvTbi0TB
Tb2AY8h1Vb+wCXzKRVOBCcvWr2PhCB++VEkao5gm3Y3ZP1q+7F9IsQrQSAly+6/Z4ntxKXzFXE6T
2aDTvyDYrDAFPBUI0SrPdA9rvepoVUAWWcUyOagN9J6OuAvg1RvqroYdj/809MCKT5/vTu9HCSt+
sYTwwjIUkU+atMNUny0+IhzuI5Pk7SbVsYKyYQ6xzaF4UZmn8YI+FtUL917m5svO+Lr5y3Xms35C
YT96/SpMLcusY0s9EE+CMGIQNgOBUkdar9T8ClbETYmh+GDMequOXcG4X/r4FIxNgzAViMHDhce9
+v5c3t4Ly1NLVZsyTnVB/f9P+VQOi5s2Mhf/0q4pdsMz2/R5R5Zg4XW46Sfj3cZVP6biUCsBGz6j
6HxnmES35AKrNknFih2cUcxBgvXtwJWgiMCsmlvGt1/0EVKi6TLhBSdTC8KNiJ8hyvwJmdBLGyrX
7s/8wKRCH1HtiHEkq2vCn45yCa7f8gSelpETYWBsgJVmSbY9mrjBn1NxcPkBQnmD63YyXq7I0cxN
wBM6mzpplv4VexNCLdDVWOLnyGuty+6obIgHHchqdDGvs2hO3q8/NGE3pi9OvlNZOdjHYdggWUZ1
ld9JfXrdLvfSGXjWDQLTENeP1X401qw4VkvyQzouBdvAJ0jCerOTfKUXzTppMM7n8yYNXYlpdE9B
a5kl0UI7YCugHqzPmE/G8VGQEPfunkhVXZBywYqBebS6FnMuMCSq15RKa5gNPC9nO3Ao9pjNijHg
eilU7V1huDaTgd212AKRBxdUrkPNGFH/MdsJcphHWERYJ+b81BCnViHoptQAuYIp2PFww6828rWK
hHJMQ0i2/5MbdoNX1e/PIN2QHd0kF5SRpqrERylcgppx1DwIoI++xC6SZHzjgB3zWkjDcr2Dsxrl
zB5YGq8cjZaRe3j9cByk9G+p7ccrVnFaoSxl0O1si53OdF6/4Iyit6rYYm++CaFRHuwoJIQRxkDp
vAafb+505QeSfhwhHrtO6RkIECvFv9Ab2/JEwanmTB9T/CG0hhKsMGrE+Qsl8jvaI7rgV6yW9y01
DlVSo5B7ea9jA1CRdc4iM6BAVuMoxtuDNSXSfYHmmtyzhVksr8lErihUEr+Q2IonSG5xbXsWquuh
EiHDKc5Xaxv+U5oqXlDuiSZfIdR6t2yyRfjpV1Sqn1y70pz/4H1+CNULlPd+FH9ACDWvpKW8ZX0n
qAAqfZ1qzWpohJ9YO3YWK/ZTaw2zgkhYfXqBgziA6zmIHtJICIFD6bYW0aOaFGW/Y3uAyScotoBl
6/DjdMHs7Tt76YT1jH+l/PUUZwn1xt8GchhMTqIIr0p8CDl5+K2/Bxd0MEY8yaqUenSXe41N2Qe+
4UlpedquxSPkTm7AhHa5lb/Ihgo4jHhQk/2krOq5esqhmo8ukigEoxsKCFEXjnwKqPxNTFkIiygY
l0q0pp3FE0mbm4f2qlqKVk4C6ctDbo4RkV5anViaSGP8QYKkch8IteBVke7HdvX8iNoV2jlDU2Cp
ANGTzPA3O6Xqj+Hm92VP3mbo3J9BGw+9+zWqIUcPZzP1vY3qH/5hnNPytuF3PWMZKhVfUSI5iPC3
ioQcA8S1f1Xoc+duO8gq+Ao+IQPZqsCJiS12hTH5bHMDprAsSQuQBA2dH+A5/LXpbFYWpLw6uSx+
vo/3Pf64wmPg1TouGNWFnLr4OZOcvKLaIYYVZyOcuAJ456VkAackYZ+bRGiHAMSlgZz5FRARJkO6
PkhM24rjtGuc+EAnSsW7d/cLos9BPhqP9WGAIg7RmpOIWv4V/wFwirGu96VvQZdcgoOFrfyWmjjc
S7QoXnywtnsXT/yLVKKhdxeKxVvILTlI1k2XYIkyw7TksikF98hhYG1tAwoRTVhXQHlN3MbZqhj3
EE4TkyfbdqQ/xG7gUyYqTWodM+AVqXhZFhGhNeQ3eOmZrME5G9NzkzcLHoO7pI093AW9gE1AiGiF
1QRXhwqquTuZASTUCUQ381xPxxG3dP5iCV0bveUefa0my56VYXzUu/z5n+E/Uxa94WyxAg4aHPtO
McvsnlOvd6l6h58AS8YDgar+fTCA6LmAgFF3shZxAq6M7lKh0DWzGd+fnW9Ez0lcRwVGOs5nAPEn
7UWKuHvu0wKb9nGQt94LN+jtvomb8c38J4ntWxUWZi7ArieNeJtIBPVgKhTFTQcDhNNURKQDU099
pG2RNubjDv8XdJocyzERs2xhNtRY0sYy7Dt+9aE9pmTCNFus+d40zHOsfyGUBRTMrNUo2NZorgrB
OFUyJdQvIaKjPMtXrgSG25eJrStDv3hnihKTHRfiX1njWZSkl4IjzZpDS27moWCDDNA2+Y2XDOaP
jfZ3ZYcXgaFU23EY0jJVRJIA0U5vcjVnJ5BKHCbichTEbL4qfn8OYpejA0LVOdw76jUTWUP62j+w
MN7a08Tj+YDnH3q03bvE7717/lGewHk39ESpLrAOJxoPhqBIGaB2o5vVd7xzM3dVVKR7IH1Om7oD
LUAaclgCGDDfYd0ZGvOqoe2/C0mq6MIoEXa2QPCjTP/eWd0N6Zd85xCUdB7ZPbf5i8XaVDxojUKm
8nuhwtZKxiKFQsrm2mKsEFhQIYy6c9dc+1TpJy5qD8dVrOATRw8MKQ+LpcDOFE/Tbzudirb1LpZz
FeIqWqWx8p0tmhk83zKmGv6nGexHBIeY38tJGhus8GfJ4DwDj4riOpn9tHkA57ad7MUSuSMGVI6U
4MeTrWazko+RrNArVUFP45PO0n3PArzlpyGRwq85eU2fkSC1W9ji+rSJBfqP6FZjpMeKyAXnFoN/
EJ/DcWAtk8gqD2b2ybV+WrHjlA5T/uuVgB61ucLbf5peqeMDIPEWaSZ12iv59fYUKFdQOoYNEeCs
hXLMu5KXs6ZDxNFhokICPgb+cv2/Lnr7P4ASbFqMoCZ/Fo+MSJC3fD6HoV9dgZM0i3z1rSsAATbM
PdkYDqYcNsvCjFeOZg9OZQXEGCl16rV0RmLPvoH73xPp9rBKc2jutsC8a8hqio+ddfIQjuVLe62F
jTrL/n+j2R6IYsZn9xjkJEJQ/aGK30ZPkUGOtkRyvY3DXNiFchCHhjNbs7QNI+PisvyeIhGz7AGA
bKXQJggjzvMxPhit6/hIldGCV/qDXoMZHlfuLdV41WrjGKK1BITt2Rfarhzo/8mZav+TLkDp03MB
HU1qs0t7h7IOhL4JzJrfBaTryT4pBrQJ9s1B0TckQ9G3Yh5F0Xeq69FrsCBugzParEHUGwiIaxvt
odFHdfg/eaNfsZNvY/Nwomv4vwc4PIuR3lvrm7ci3F3k4NjI1Vh5wCg7mD00YRYa73WwCs6SGCeX
Uxm8ES6qWazN2+KSb96mkkh5KKhCeJKaqxbFQAZg0BmbkQ0b2eK8CtM6Hyqjse7jzZHwo+m+uXnZ
5ClD24GvFY1/NlGAH5nydI1DvnIvyyoDrTRqk7SI/vQO+A/JHQVZnnn+Hph0/C5412HnxyYeQa3e
ym4lTBRUcEV8jXbz8bYeA/lewJYP2jeuGv5nmoQG+/cXmHTM6WmxttYVdNzzapySmSwyvsidbVni
mGI0oWUf+jOVJSNSGrHN1Dv6BshOL4/B+znslSywEONrJBZv6B/RnSXTd/gdjmYaL2TjzPweW57S
y3U3YatXF2gorXRShfbVJ+SgtFTReIzMSTwTgUmqvma0G2wQiUN/emj27yxtCs6K07nk/4gbe63t
JW2M/mx2PiXC3teF43SuGCg99sCb+WlwkVQ0yZlh0QGSuojPArp4i9FgtY7VzNXnUveceWDVYUF8
S9j4jso57hV/8As1yKECeT0IH6vQGyxGNVfWYOwxdl8+x1vm6s3YNHpTrAJONuprNfY0bqaxDuDQ
GYjciSj5+ktyyMxArdVQs4BwV7LPY+vxpik9kPMOe5U7QzVzQt3nEedi5q29Wnyb5E8OPhQhMhdX
JyCkYFWn4kFSXJLnealkSRgnAG6rll7DgTl8QweDWWg6iKUERwIjRAO6COixWFGXsx5qlu2C66Gf
u6BrT2pLxYe5IEM4IJFEriyAV1yCQhnP/ndDp1CRF7U6peMuhC652YDSJ3P/dnwjFU8VD1dEPbol
SspunxN102aDP2tqOnfhlJ2j5FiTGb0Mp/j3fUcD5BYrW3U+gdFBRy+xFUN5zoBGQNqkN1yziKWi
MMHLTsbV9sY7Ci0abkkIiPQn9h0X36wVncFBORgsdRcnOns5vdbdNj8u5c1teECNDWKW5UJYyBqC
nPF88+JTpE1IgfRnGqMxLlKnY9wzUfwbULe/CxB8lOhVHuUhlU8D2+WGpA9STOjryTicaeusYnzc
996ZkfiTyg8dX9VR9MVrfhhRKcAy+/KYKIyJAvgdJrVVKwZYx3GB1Gg+KdG0LWS3Fp6m74qb1rcl
pK+Ll2vJX998GeWPP5jHwZyWpPF8Yt8io3bVUBN01OuT4TEFR0jEsX8x7q422a7yX3cKmFxn6B3P
32G/bojIUMSx7nRYJ0usiSECh9Lmbb1EDVluvoNbvxDt67wfvEU6uxF/b5zILVupxeLRL8k+VzuJ
+nY89KUQTv6LFE2cKq5IMaPq3JPRy4iv95yzz7hIv07i/dO3oFriaIaxZwC2zoBMfDn8qDxcc0jd
cwLUdIJpQ8vBBWG97XRFgl9ECXkNDR1vNzmBnhwiAa1OHKq9AtEJ7Nl1i7Un5Mg8HJtXkFeNnoju
kjKuDupGpeZL9ag04sfRGwh/L/Zw4NSS0AhDXFh8SSgs7uYbLgMC1kMjrGDC9lL1y9P3zb6vgtL3
xvrRMQt2f2F7Z8X4Hp9/DplrT0TMo912ZwtsdTNea1sTAPQsW8lWUlChsffTOOVpX/cOKFdvV5k7
9JFw2Br1fAlxxVKR+v8M2MflFfBX6/CQT08xKee5s/4dd05MPlMmjbP7lM3ZyJIbrYDtgoUwrhzS
WHWnh5gHi9DaX2iNxJSFC7BzPVxZf3vMMg34DdM/r/cJwpfX/I6JaLfyP0fgX8vLpJIAUysAXkuV
c70/if8m9fSmrnYrsXUUX3rtz8V5B/83fprX6BfSq5HrSagPzQwqDhZ5ShuZV0l3rB8+5sLD3/oP
Yhb8WO6axLb7YISUIo4NuxP/xcLwiEa0GqeANt9fqYxJSRGWlnkQC24Hwd4Rz1v5709FSlPssn8g
18BZ2fr543f2GQMDxJnH162m2reZVkW8F9FKJ9oLKPCoFfAOKSALtF24PPGcVnHLAhtx6W0hEbSf
WtoyZqqnKTaZ9ShYOV/+pL4GmgGdqp5dnalgx76YDIAQHAG2eTWXjbiWCJfmr3xWY5fXep9fq7bR
8sSKeiHaIHDXHsQ77KhWDfSMjW5tCMeSXZCYjYNcso4WmIno6qELjvtm55JFiYyFlwUtnEIjoStB
XLAy+OYoCF8dJ0mST8v9dhhHbNWtWbmR31S65gAldRRDPz0JswFZS7tyjL7KpM1/I+vf8JkUXICH
ywD7iLVP+H8/eGQ5C2PtXH/lrOP0gIE9yzr4sO59ERhL3bvKhgU/nQs0yHfMChd4vVrzbfyRcj2g
ichCsf/bJxA+eNrwGOoS8YKz2Bqvjgirbub2eJ+/N8XQ2w4PKaq53mzgdcQesOr+H3ubCDfoBDIl
n+e+znP0RREHgEhKpRZ7H04bt7BgyHYqHyqKTFKfi/DTxBQsm/HlAqEFYgoG0KRjbce6gm/687j1
UD2fJYYhMqL5QF6BuXTKw0M6JcLolaRsd0AeU1RiwcZ3H/ELwy8mRgJ8uBFr5P6SbCwlG/dn8rUb
0IOBV+8pyU6o7ByvO26BeSLNH6+c4VtHNHn0taUgh/t+X5fgtAbSHzAnvol7lG5VCBrst50GHHII
FqzaSjPoDRplosNkjh4Oq1YG2w/kdmMFje41ySar2UzuG4RKpnfe3BkIJw30d1qIGhiGoHR//qs3
oQVxLPta9FRHqTl7tCDmTjTtEkH0P1PnTRWlsqxGJ1017IwxkH6A35yrucAi+SpPJB8TX/QkwgxQ
oiOOpk/aTjyduQhIksAOuMxvHnvZ45wrGMor1y3kphpfbsqxSMnP5FO6wjwqLRnh29or/JDQRohU
ej1svNWgMJavmxPcnntaTGWL4mSRjo4+XkMYcnvOSpIWOn+aRO8o8YLxNqsWlJ9fkaZr3dV3VT9n
I6VVRcXUkMOL7u5QMZ8NglcwUahyalA2vXmYCgQ3J47+DaJo8hq40qq4beyHcTAGDYCYpomAJk+l
gF+GUOjOwmjDjQzFERqRu7iYq7JdjpWqckAYjkpD67ueY7i2l80I2cQAqckEH0fk/lv0gSlSaJQw
VsAObbDrKTeC68mdZnbN+LbTVY8WxR33ekQl0EV6860/Xor6EzJNQuFkoaFkEmYUlhT19Y3FfCy6
CL7mPgtsDG20zhHJCTObV3hTP5yVqfZ4289cy9xyUPiOIbNDoTHqDml4E1rwTB6P/vcqtiUboFq5
xUuD0xTWhva3XFVkwwZYX1DpYN9g6qU8MdnUL0LIyNbJmtibK8UQD44U8A7jbrj+bndolf7P8O5H
SMmayqYRRdwgpRMOYvospscGPX3N5V6mobMqmoQiS1BfbWqA76AXr/ntKxVJSwIZByWXH86+X+6y
wgYX0Ol0LkHVf/YNdeZ8leKeW/vx+tU2NTRBMaSHo94nHoOQ1RdKrZt1oUyWX5OdBojEyqOBYeHT
YWwNniCuRoIm2uIVcyuNQr3qQxrWZdnsSGlpRFOx3mE8gYI1p750C/N/MNi4oD/dr1e/ZKhUEMyk
Z520KuJXQzTxiF3f9aQMKkGc5FcOXiJQESm7iTLNZleCDGsFolrvHfyaqz74HxnHCMDxfpmD8KbV
ks5Q+f8WstPSCSv+JA/LOJlFJzNH5BSf+7nNvJdWCn2Ti6YojjM9ehXZxqJGk/rnYuVGit0K7bhA
SvT64zxZww56Y1neun4zZD3/cuwp5fiH39sMBnjZ9OTiCAvaUZ3KlYHnqUXKen7FPb69bXYaVGa9
QOMIkk6GRBRBMfoVQNMH/M8HkkRTOPbEsJ+q4c/uCB9miXzPPYxtdedEEOACWz+69bomh1zgq2jV
Hk5966BSTRnbxqMnR6v5ZJbYYPNgLTVjR0AptAntnGIaaVD2Q1kHf3rkUoozz5dYkLR5JZJVLnb4
EmZTeR3Mm1X+uVmzE/g/izj+ZZaLtDlgNvIrO9ZMIpgeq3sr27ak0+nzDJeYpHcAqWT2Hd8RxH0A
W7/Hz2kcwLSs8WZw76CS09+daXg2Db3P30qJmq1DkQeef6MRHPWnYgNqykG+EJxtYp/ympDBE6pX
PpCNtzXT4UpVoAX/VO2eBMyRdId6UceluEDcrHp/cCaDIhLlN3ULkuLVTSRucdY/hxXX5SwG8IYm
8WTOI8/3QwtvKsWjiTzU+t8UpOAGkwa1CihyrL5WBkOJKrb6wm93UkkDd1o6EOQxz12NRTDmUnLo
nM0dAVchV1FixJvx7f72kw9w3yIDN94f5EktOnlBrPQOVizfCBiWUSO9i9gcBoeT+VEsdTM+FIRh
zWjmiuPmuu6qlwsStxXc1F4JJEuowJT+4ApFVUO/3MUfHcJXFj+7zDjmKJxjVO7GZS8wUfrdE4TL
q5vN7rlHC6zA7qfQOM1bSsuZD57CbPG7KembtI3n7TjGvlQUBZbZkHwFxgiaAdTQTyemEkWiW8Ab
K9saRBOdwqym8WMjEp+cmg/ZlTpF7bRfFySGfw+cd91IclJtpappQHfizxQNJrQMfuUyP4GwrfJ7
DNjzO8h8h5OOOQAo6hmev7N0q5jdLkDTxMmasUz6He2j7UrKdWl0jJ+Gx0OhHJVIN0Whis9Glu8y
wcU6N51IaAX0cC8aHtG4GwcmhoUQhHHoJel+51wWjmWF4P6yWjMYpTeVVIRHDg4bFRUFqgCkrusp
tYWKWVNK0A66qbV6j/QkEg7TNLewCXCXmEmro6hadtbmRZ47SXZypZXnC9Mdjz2nOfxpjxmfAWwM
dkMtioLDb0kEQI9ve8+KH0B6LCBS/WPFlsZhxa5fPROdZ4c84yTbFIXRkv3gH0jCoIixYyiTxg+J
7Pu2MbvsFlYQXAvVWOAZ56mniZxWIoDlZycBKzrt3y64jaI0cAwsYxVnSSG/vDy5FCx51kcg0BZe
RfrEqr7Ul+3la1u5c9jvN83+sVepKXNGDv9SzWnigusffqC/f5GM+9f9Pb/Cdj7HvbKLwB3AokMy
yopbaZOX/yWo0CY8hdsU8MgjfLw++P+RyrNFh/58sQ+o5gj0r0X7e78EX3hRWFt1TQG6HKfUVAe2
p8YoLVQlzoJ344VA9euzjGS1ODptcPUTq22u9cmtxYz60ToPDynX08ycaqwbBHAb1tVpJjYvH94b
1bdtyhKx5TTG2ebzvemj/g7V/fOda9rV8NguwfSdZivPGs5cCqBOJHXlplMrnwCEYdrc10Bstk+A
4QKL4F3nNFxfW4wimAnUjpS+ashF43AE6UPeqFlmb/Em84TexMdkpqgYXiFj5E3u2n2Ec5S2bqCR
GkoO1vJJvC/Qjp0mffy2v6puNJ6p8smEuOedBRYteQjC1yHyMJFV/+HyuAeaPP0OABKDzG28BsEp
mxt801GTjxPcMhCnUGIchjXa3HR8YrZl6BQOEcupPjpM3puvbLNDRb+P2Ylac1/BB1QUgqD+Ak2e
J1pR4xgcbfC/uFtRkd8xpv9IKRCYRg0nz2HmDvF9Mc4oKT4zCadb0sU/4lO3hhYGODYH1d0HgcAH
L5QhXYGrP5KeYNVqWEuuUsQ7ncbXaidmCyDsaXfCpRLy6/Mrc/rVK4TltOTrNr0S3AANT8xzdUfw
4rsQPI+tFqV57bWL0iLYLn4Yw44vbHybNw8UpP20T6wY3yIsP0TYSpfCElw0IYMGCZ4G5izvOnyD
Aq9t/9N+pP/ctrn3YBSv3Yk0dzDRwSqUf6ygn7zrsXtkA2dBCV9I3c8VhNRRkHkrpToYJjvZv2Y0
zntAqU+KvfD3ctZafECbw2eHsa2Nm4mfkIfrMXQCqmFoTX/O9Sj3zECoBOJ9uRvgWS5dfPrmVdkw
Np6An7tic2RhW32xRzv92CZFOJ/aDwFy4VITEO7lRfI7zFEwT+KPYybvaPqpBzmsBY/fOeFjZfy8
THLoduBDJEOPtTZ1un1cCetgMOMouhlBllT268MabQXiwghJaRNPdr+6JrbIk2bRRcHOBitKKcTH
cBNn/qIOF9lJjFy4O+pQ15qB8uHNdT6QyffjwK0uMHJIsfGQRh7nN2/Yg5aXPWvgAYxn/n8xhP5U
sWpSl4hsa6zbRSkwrQTSXR5MAWehEHg9OcEGvudduzPxvV0x8pO+iDmsD1EnRe+L1HkI32WC36yC
s+v1bjR8N9Vf/UJpqOwPRt+JrgSGRGxeCmZgPdJFlF2gecslOJFUkm4fYuhR7dIJkDv/LKBuwYJW
TUJXOhyP7YAtdzMtBKskZQS6L38Xx4x4hqYEyX4pO3dMxr908ICbPc1KrJ7FCGwh7CC/FEQBrij2
6LbyAJvdmy8IAZFoUYH1/sKGcHvsvfLe3JA70PtyOILx8OzIIDBzbD2IuRI/V0zwnd9dda4+zcCt
U77qP7+hg/qRo+0/3ZuDo2Oz+U6BUoP2jqRmjAv0KkXf90nrNj4m5Z+m8gWvijuZnZKRkGwi+fb3
0LWMFBiHJvWtfP44y6e99wvVksWaZ/xE9idm8nxuGIqkp4fCB7+r5OT6heVSWSFuZOTCzSUL6YYG
jsoJzxtuRmRGHlXnXL8qbQW0sMgS5yrqNcQjILb3JPeYVUhrbAuwhSV4qEWe1bjz2Hpu/Ai2kvBo
hPnbaxXmGaPZHw+rLrcMha73HXYAmc3e22AXh1yFyNhHmR4xI8jZd8c2F4h9gelR51f8ijXFzyA4
j3MGfeY9O3EZiuA4OBLZKuH2notazKWVlbny8+tl2DMFubha2469rLOfeaxpHVO3KP1HrOpCV3hN
rj0OVvXdI1emDYSGCUB8QvW/Q/u1S4PXMeyZHIqW/QBDpUfPWDj9QY5yE4JfKRhDRfM8QUXpEoRd
fhEovoDBhkdA1iM3L2G943K0paCNgcglXDYD6ykYebpdGB6aIPOhJ9tRLKg8C/Tcd0p0y9k9iKC3
NaVTru4peVmo0i2uChyg/vvNoSSsKYyo2DTrIXdGLwum1dCwVnUNQ/TJ2oPiNSUnH5k2TUdz5ryY
6yJBGygk6y/BtplugEKMEurEfwlQUAs+aeTX0WFZcY8NcahPqeCv1La93XWeSf31UthxVvd5xvjs
htohTLT1nwy/UDtqh4Q9GzweZlsjSO2PW/LG6zaV0xv98/iHAgzom4iU3kTbrcbgvllwGtBiO5U7
aQYHV5C4Vfwol+esSYL8X7Za0R8fbD2/+EJIm1YJH1YazOiDOdqosr8/KBR73w1V9frDqt01SWui
5rAaKPcAYDFyEM4c+/BOIGYm+FKSeTSsqzgH7zNzOcTuGlcJAshcoPllqUu877cATp2XbV6sF+nM
kiIVd9iBzmfmTgVBkfU1fdFyCwYHd/FdsIFomIl5b6YfhiCm3KnM/GDrYRYjx9INYtdMEK7KJfmG
GIj8KscViQqDB3sPEu3fk1+L76sR/utazSKz0KpIuNYoNkBopqKJbeHyE9+5+jzaBhA7yLLGADUQ
jyizQxLRVeemLNg65ALW0vYuimC/Zc4NShYxr/ATe4xC0wLX7rOLd13UQfKtQZzx7OB8G4r70seJ
EQcfxHV/xp9g89hrQzvFUeKCC6ckYxl51tTec5K5IbhIrwV8JqwxIRNMpEGdiSon4DXf5fkZkJFk
ScFQS0B7/rqtezacZIMl3tdFIA1p9/mqRQepX/Ei3Nxo0KrDghBBQ+8xDWYprgS4jj0W689X4PMW
swEEUx7sHwsd0PVNIts/fm4IQcRNL7Rf14nO3QSc8590fU+tf/6WspK6X/zzdghx6AxINGSblyUO
87pxcnGnI+bMDLm22ITG1rgY72ouzqjLaJa/6uUYu83dttKVQrOLzXi62Qqzz7YsR5PTMIPFUztP
/O1s2JUvHOl1d+QkgZ6KcpsqscotdA8NOKWsQrzRXqbX1PEqvEVN2TYUzEpnIJDFvB4EmJM/bpPa
SFb/SCWY8E/LpucWK6PJeMGE0Zic4VShmGBU9FcNSJcrqfUHZbJivF27yVyLrKpOm/pZ1yZMex8a
H5yJ6+Gez7tEnPLl/Br1ua152+Uc/lG2ESda8lCzZ9fhrhNrAT00mMDVzJGoV9YuQxjXGNqm2KFE
oaeDj20A0byqHf3k0dvdEqn21wq52SqGTCWiueNDLF/rxBeMh6pMiHQLhRiE7GOeTtVNgtaEH80z
e9+i/+38w7dLtvU6LQFTyUiy0wkkjrPihntRoHXV8w3L8D2t4Hy0i2esa10aOxHeoxCZy7wi95IJ
r+Cr094QRqiqhqT2RkMoxcztUBMX/txZusISwbw+e8Ia26w/hERbq+9mbqKq4Q4vhpEC2n/XI7LI
O4nqUyKX4sqcE2oKQBaRke7vSdFpEPKmXBjpruUF8/FziYm8shG3SjmOzPB7uKKIglOhNXqHA5HL
Jy3Lvd7N95zD9WWmVL6lxqWCGlQ2m3qfWdaRmpF6DzjKovVa1buCx4PxRw7gdsXU8fOEFg+Ol7mQ
2FjOXrpby27K2+svd0WJCVGa6kQkv1zduN9LfDdTrzWtkZMUDG9TV0eVSiWMTV7mjJpA2jUr9q/+
66Hrn2wmBHMGEJNVMSoSOqOY3gpMFVGrd2GewC8BVEHVJtZbTU6sFaKZVbvixcZlEBr7STGETrP9
hMI3g3LEtgTFLvM1HfSEs9rm1yY4yhPFLkcUp5B5o1zxh3vIFLO5ghAPGvN83y0wpcxfU3XEA2FE
PSMBK18/pIiEVHzHgCtrh95SCuvcWAhVB9Iv1QxEeVA+w/1sko4xER5eVj2EBXyU2v4FnogCZ4uM
1RmwEZp+dxbgY3P7k7wKTzh6XLFvH2OQudJiTiGvLMMYeyVwP/aOrzWpnrVQTbn32mD05Bs6IOLA
ibU2ayQVLmYFXxwF+UNLL10tcbtyPWnIJh4CbGXYosNaY3laG6pErQmfz69cxNugqLtJX9xEAkao
pbhOHXlpL4xm50PN3PJpEwiXcnH51AaVnhbN2w2WDWIJD+PWnwQ3m+/eD1KIMurpHMVDChrFTlBT
ZnetTpDoSwSIcYM744Doan6d4wfpSinDO8JP3Ucp1a4QGF/ZqVPn19FDRbAZu5fmxd00rLbLakkx
iIUNFmgnPBFx7Yubiao21+M5Kribhv1CjU7aNcuNk/Lev6uiciy+wEh3khtft2W/OSuc0s1bTL73
xPA1ocgjs0pb+KSsC8fjyRFKwFga9pQR13ZnoWOvU4edg7m1BxsdeXqcDwD3kcm3m+Fxf+h+Y7nU
MXPlhvMX0vOLQoYhRJPKlY6yyptvQ+1JBPzv948Vd+V8IQaNCjDZ/UlJXp6uvNPM4BLWiO3/kJWf
ged+VrIdTyLEablX9xuxT9pxd8aXWU8hQsb8ERH1BofMpRWSfKTJUhgcMIsTk5C5JhfQCQgaOPS8
Sza4vSX15TjIh8TXHIVsj3/G8/BoC6oJvfFucxPuXiQlkef6dAtPRE5dPolBDBF780kXYdN6gptn
XNR/zhma2uA/I9LmWIMn/ZAjDwuc2n4dyCfpy5YJaeVkEHusU5WrRJxSy5BzAGKfiTs/V59lv447
QA3UPAgfq4TdKH9zc872E1GGCdgT6hPGSLCM+wMfje6WRHogEr+nEzDOlxw249tgLf/t7qlzQ381
AQVt9qgyMKw6Dn9pb11t0N7zxi+CJYgTyXjNOKV4jfBfYS9WQRswP9w6qIQrX4efwclmqngm8hVP
lIwKvwpkMw9g1lbAq92qb85AL5vNXNCHedcmIU48gov9LGtvmF4nSYre61E60656wwMwq+SMMYok
ZesRmk5ff5/AoOlKA0Dfwp7V2FDjTM0fQ2QbrWMTsjwQIxF9TKeMkz6rHEBsqAyChdTviNHQNX2A
wmLFxW8pfn0EwN2ChyIn+cB5LaUMQlAYtBP3kd/MqPVnKgG+oqYr4Zmpv8GWMF4IFvqjTmaWyK8u
5wMaMpFFTl1siQizEr7gHoWtucs13nkstBdbyukfHyuC3xwbCg0PAaqy8UlF+Vk1OFt08N25fBLs
IEJsiFJCzZGQ7gASVuF8gdyyP7WxK2+k8B8sb/0bbpdthwbFRmgPs9iDBNboEq0L9tisax240Cu+
F9ONs/cd2wuxkL4pCbCdK1Aq7fwkHnLZQ4QRvrAACYllfavBSaPLmlVgIycbmx8IKsUyA0kBnGlP
uer8zOP2chgEnDfQRtfzz7nyrd9JgVdjwFfUNXwR2xYOuTk11qy5m4qY4mausRneWidJnNRHT4/T
iTeTFSCG3JUj89BerU2D4IHpxeXXSVvVyTkizlOTmBEH3alg/54lS2uoMr6XMY+VdgtFc5zTrcZW
bwb2KIZchzrv6DARs4Er/fun1vFurT4X+0NkUnfTOnM8Ssd2qOtikXOI4/VONUc2hgIMEf6EyrZO
FuuFTKQFSc0YNHs4mvQXqWGVi7lRqWMmSZc9rJkZQXDuiTb2QH7BKRWfyXPS0YwPVouCY50hEZiz
5FHkgeQ4LvrHHyKDEDPKeWWheM6ioEhEHJOPxAPOFeNltQv54KHsmhqvKKhTF5/pJpFEzpMsdDws
/rkVwT1eWoAgvAMVwcAuS68nmZgSo5+/X3Au0b1KYKtuE+7daqn1ilkYKZ4EoJAx1V9gx2Ehg/L8
PyDGYPjNElx/+ehe5pRdzKyMlGXi+/K9LuKMRdORHYHB/5dYIUtYnY0eKfpb64cAxA8o25sIMHRW
qnUxNuQj8IQ1aFkCY7CPTfw2rD2hc+mrPL4w36Je9/JU+BFDbBBLLx+3ILytMjbnBlnycQeQNhMC
Vk6a31p4UILnHpXWEBR6PqdaRj1OAzxl/kGwEgkJj/nmayjDyJQ2CYUMC+aLBhhlYLgoeDJVXa5Y
qDDRsDxETCrDIRW2eJDYEXyQICpyx0jQ5DT4ZlL4GtGFyWWbR92tdPPcEByHvlw7ZXATjmtmwCfZ
r2BNe8B3rL/+K6ghGu3l09FcZRifCJZQCX86Py39tEjwAkvLo01TONtfmseKwtGYP4NFjN5aUO06
5lCGj8CtZJGwjoRGkiaMN9TsmuhmAnbyw5cIfzBhN1GLCtbZB6fqnIXL+T0wkUp/hxn7QUpiNIR1
kaj35yQ0B+D54XfHZS6xjULZTUGxxqnFlzevSMvMh4zNXh1OyjooeDoVxWndmFI621H9zDx2e3Vc
7z8slkcbGIKAipDS1LUkU7nAklqSjg/P4lMgAD34Dp7RAjQIyLpL2tsJ6khO5tWGiQ8WcFa+iF59
Q1Tu/50eqXSFdAF+Q1LnuZgpnKoKBjz2yqwvxoCUPb9e+LdVhL7oPcadiS3hapT/dUY3b7do+Fe/
Y8YID/Om+zOJM2LQPPjJAls0ZgSo/Czc4rtD4AFwBccTbdH8ApGZnBtpoC7Uk0AuWwFlD6j7vgIz
DkrXNbe0L+guZdQg9QT5WT9eFRUFOChcO8eyX/BHlHC9PE+4iLo0VGm1QaAmePuj3i0C+wxptvaL
ihyL8XIadp6L/T8TKJXUCPu7macAJ2ZCvGBAM8dVAezYtbFxX3G02Sr60U80mC1kBZ4duVu8N0T3
zBb99x1WJm/RknKpV1iFqMAwzyEm7vy4GcVq6udcCLn+8MycmUmpfIFu4zdks5CjjEdA/efxjUep
WDkVo5W91fAY7uxoBQN3k08JHRLhkCpeacbF+ijsh7BK+6hEuSo8ENKx/ehVULCMn4UBUqkzqaEV
P8fxVjIYBaJXhHuCSYX+3p9iA2egSUMpa7o5vyQpMqfmB5/duheHJ8Dr1CkveGB6OqqM5akxUBRa
msaP9OrIlQ2DAK217dii3Tj0e31NPc2T/1nFrmlFMm+SxrciLg/He1yHK9aB07bvxV2w5x5R4zKf
GfPFraBDB7N6OV/MPdADiENAnX7CYKjTXGov5M2OYPqvmaMsJLzNDZO4Mr7MBcpT4zwvw74lodYX
PhKFCFHYFPfb91mGNk9WvEPH2eh6EGZAYfeRtxDYCC4EIlxKi4QkHGX2EDIMWTp5q60u+4O8Q4lU
mUDdA65THy+EvryJBvnEkC8ftaABrErZtXctdLOaKatAHvnMo8t8G9Bp0DxMrh0WppkuUCzf4Rtp
tekaxUVbNp8naWQWus9xWb4sefRodnGKaSgNorXgzwi9hz/SXCAGKwig+bG2DFbTlo8+gK3+C2cL
R9PoBTR30MaEFgGVD/ylq21urzABvOtt4IhSqRNF3m6hiUzGdozSlBQ+ADGF1DQnoYCFNnhbU8c1
9rvKtPfFUcYIk/EsISxlLVs+dWCMJtKQ+vMsTNIDsZu47VchThg/Cb5BzqBU0CLxh8vuubl/4MzA
Icuf7xUGn1eHLP3stEyCK721UCGJFhivzUnH/c+AurNRaqBroaMAd0aVcRRzoiFVQ5LEuPOXijc0
O9GFbP8+M9pa24a4Cws4lNcJtXq+ux+dOI9obf3yCDfobHXfyrM4gZMcVZi4dO6YRntuwRvX8F+N
aK2maS8YYnyWDGwzUvgCkJFLoQI03CqQzu07AQGpd84UvjAf+WzU/6448HLKjN7uaN2PYuWNmtHF
l5HLXayM+sDb2USNHbrziOXp5Dspyn4oQgp+9MzUzsdClhyYPfqNw2vWw4H9ofNgya3oY9P/PO27
na2qmCS7n6/g0Jj4wRL42CsTq8mDVKFRT5Wzs4WnyxhX0cW6BzU3P/SJ9M0zrCBn2+R417IZhGNi
yv8ZgSg4m+/TSv7WCaKzbRA+LwVh7pVvSSM+fImDj8OKGpSXh9ANQOEhBKNk8reWl+z7jBlYJrPq
a02XRB9e8D2UiO0eugjAU8CedrDJGqbsihaBHYo7rrlkM7F8ze3r38/MQ0cvlioF/jHr5NRQ8ftb
rpGMPt/TtXVMdu3TzHEn0Rp7LSwJBGgJQfWfGv5K090LJ0FOM2Yv28JFIECyWF96RYSqNdceaVgL
3Hbb2S/IkbrUFXhheh7qC5LROkve2V/AhInaUt69FJ9OPmPhVYunO7LC+whDEqIRttzC+lCmFRCW
m5Il/It8wmVt1RgRW9N94hLui2HdjWj0eT4EYz8kerTjsAKH8o2qbvjDSxfgH0YtvJq37RBQnxvm
8N+dGvCNs0gPwJ6mTVnpbUbty//sBLslC87Hb5LBO1sl7noB385kB2WkjmRmFglrE3WG66OQewZf
rSvkK14CWLQY36oWHTj7DQ4NXwYE48ZpClbPyf6kl9HPcBnkYQbNuxkiNJXcDzLIvlCLcsD3by4y
16FSLR/VrsE3+5DtmBwQstzE3lgBvJCNfpeLteljNNvwNWzeFMJ88e9JW4zx4TyVt53zKJDFAKJz
8rBV1FkcCVKUk33Qyck95rUsts16FaB/g9hJqESjWVlNMw3saskPLBu7Lqoucmh/Hu4gyMyE2b8g
JtjPm3ax8uBMpXkICtgqYkuZlnvoLWjrwTpVSjPreiY71A4Sb/Qa6CVa078vnhDk7Bo5Y9ZYwIkt
j1NJdGctLdKxZP+ZB27yKFOBaNtmPaX4O48SimvqUMTDMK26sXUGpAh9gTOtKXnMuCTMLutHLxl6
C6jRg7Y2QTUTyznovlyN5OEYOqFbgFPBz1lxgMlborGTeGiHNArrQGy/rT8GPXl720wHDIpP8n8c
Jw+Cex8fj+SMxtWqYdyaUbp17GZ2uD8FiEnsom9w0NcCuro12YSwT6wagTmHvx/u8bJOROVa4yIe
83vQ6M7WAquXlNHjCRtu54IcO0vRMqBbwJUzV1ega0gbtKY5/Hbmk3LteD/brF/n1qUsOVxhGeoC
zsasIrd7xJo0Wj8m15lykL3r6Z3OCBvjJdOngyWvUVu4mVCSD72gmWtT8Q04KpsPfDfrviwvzOFN
cgmwbbvawCFtBwvkC3TAEyhXM9cF8AS9BxaWw/WuRwGNMLDLVsJUd9TDdgb3VtmdKbonSImKFmy8
S3fzpaxHEmkyPdR0e/xhw2xLTg35Y+2EuEt1Txq7Oqk2xCIt2NRff4GS7taOyhLzZ+hTVrFJ2Sva
CnBdYWuObdIcQ2ipCER14oRA+csf6wti+vVzIcy0etBkJfre0URFRXlKl5ndrNEfMzxsH6hQelO2
uSYRs1sc2fy9nd2WFbO5TLyIKphSm0y4xXbGZ0G4GeX8qHozAfRF6ULMUAs3T2o/0KQFWaUvCUyv
3z5GBUcY+9fW9rBmV8RGo9YaOPWroE6gR1x33TUc/1UqPrDEBLUTVFomgYJBR9gME9PBTQdR+OYO
1Nj2/7NjFi4tBbA+Ju8IcJDzkPxcd1YPhLECleZAFXiWk5XuyA0CFuhkR65SjzHI0A4QB4Kjg2ZU
qs+aiaMQ9RQrS5AISxUde2xUEaL9bmveW99cs3cNPqijh4JsAcZB3jlrs907XmKce7dad1pdka+e
7VVQ0Iqcnphikym+R7c12YBIbvGG8eFtxUBb8jdGOY4qLjzJRVt+2Vls3a5AeJ1H7tcixnlB95xm
mS4Lb0zbDrFr458FJLBcppG7OXl4cEraqZtaJiv2RyLgIARtxFubpAegnhzTBVhuycPQRK7CowMz
ycv8QLb+ZUu44QbcShDw/83u/9qjsgKD7KVZfTyDWrUvLBw/fWeFqV6mZZQaF4nCTVWyQxIYzBe3
VVuk4H3x0e2/el2dDmO0SraYxS4pfHe1B4QambfztWYNQYVpsEYgDFP8IRcBwh4ddXfKXdOIYSX2
3ou5D88wvV2+dvjjotC+27TOs3ZY0WxycFTexlMFCFMXrjc9mqMoTm3MCHqtKA1cn98i5+tCq+PL
yI5RRYRjGE+xNQdmXmgzCjnahLqUMVqvSkxR5jQj1buPJf4iTJCjH0SzznPJEYmCq4ty1VRNH8jo
xguySqPckKuf0Qsb0vcAYWhGwoN6638KsKpqC894Ay8N1jdeUSbjHfBB8TsuMPQJFGAaiRdu6W+c
Ss03YaItzbMpV2KTciuM4VYgauq0txar58HjIgSmkZejI25mj3+mC+uHWSXXlYwArsZb0gdjXiB+
s4j5tjrGUUr8CFCn8HoFVHm8zMdQvUr5FZ6pqE8Oq4pQC8F0G2j5qkg9AD/JH7s9vHAzjyl+zEK4
F9rgOw9b2B37snRnWpJY9luhaL3w+mT8MwraPqBOEE5nJNaUpbkA38dLTR4T6mLUiKzEiwMPgtjX
hKj8byCLUmj4DwXJH/ZkPdg24YDTxX/9qeXfM/nQyJPdSV33ETEmeU/YowFfQ+lSs8Rfj/J1/pGC
5O0Oq03eSxN61ZzUmerF1ASgohRkiIH17s6gC248nLEEE7FjN2REMdla1JtQmLJ2NjWP6lC+bg+l
PkKgFFn44rYYBOUY3dleOAQ8qnscT1ZfEO3D+GkKPJfU0fGTIXRa5LexQOqEVDN7utkTN2zc0Gir
KWARdQID16vLGTNpKjkcxd8Ee1Ixhp3EIN8Ql6bfHqf0LCMtCI2ZfPPtDxkjDN66QL7ehj3g31EI
JV2ElQtEvPJqafdMx31RvUMq3Kg+Z1q96gTm18cvOYDx5D1FK8qmpuoczDGuJTu90gkuvMFaaEYG
g7bjwMGhk+wO2vU/js8HX3jFWDnhv9iQT1zYknICdckgXShtxxLFfVhpxP3jNgqmKawY5QH4MtE8
1gpkinYsD0lZoVUBah+z2XatP09JPwfxCVao3vjPQJTWc2nmMRjoW/9zpOkGqc8qXfcCssxHAp4K
VsJNPPFFhXGEIwfMsIpGDJWprkSmhP9ItUh9knF/NutiY36G0Ra/C3JEH6VbuOnP5hX65CwljU7D
IVL152Y+GIFjm5S42H+WWGjgovns6z8Kw0IvbkfSR6KL3DH5m4NAFEuzVKB7UNnwzdHLmAsYvY6l
9f2y9oHwNVNMHgW+lKGqzENd8nMT5zYb/smx5jZVCN4rUHYTYq/fgRQcsBwUqdr/ed/ZvDlCDNQ/
3hIu8/99uP3QSjGGwDTTagpyDjM0nJ3lbU+GtMp9LLWhWxPsHQ0TPv8PDPPuDMJYhvkQm4ztWleT
dzDzB84nynNNLAEx6cudrEcBT7ne04yEyHxIEaMj6IQAKwm9inzdeSo3p78opzndWSJOSbi6vBAp
ZIxT6lA1mWeXd40F9JNXIpmyM1GzObydKuY4jElGT66gQaDXHlwc33BVhIv32MM/vyG3cjW02lcJ
d3euwMCaAd3sPGXZCF79ZAE/U/+V7Y8OFIY/m3fVypLcRd4eluuJLtTjeYzAC+WDDBXofJs3p2Vm
PDfa0LwLWiqf5d+mXCzaA1XHxsHUmU5RqboR+14yAMdb/qBBInSHv+BOunznlSZ2TqEIphWLnVXv
QXIW5s2U86OhI5Gb6s7Yx2U3OxA1Dy4NkzHQNlYUtpMl+OKvDOPBg9PrH4sKvhv208I6nENR97+Q
r0ioqofOkGKI+t5VFfYm62Y1S9ioykQlelLJ+oOfwndydaHeo47sF8OT5xuKlQVcvVotTBygtJZM
8tMXXLEZp2wYBgTYgMQdTR43caTiaiTeiMEjAAk/IEAXvpNLZgHoFho86Y1lJPG3S6y68LaSKxMT
hOgU+17f6N3m+y9BLBFyBti+qXkITpOLT5D236BPi2QKcpt/5EW3sZ+Tcuy/+aLkMuW+eaRC5hEE
FrwMs8yd6Pn05aIONZnkZ8SL5CbEoF46x0ibk2pp6/Soznfmd9OtAXZwHROB2zqys5EforBEyM6p
LSIAm9IqZm3nEpELD9Ud2+ilDqmLoDiHoI4hhN0VN1r98wJcx+IPxooK6aDqyfgW97WLOnR4+EUC
YnqgY/RpVmg0obGfrwIFs2z7h6Bq8LDvUVpTsm7+ZPdT9ibFgtPdVhXgmieoRxJMfV9HIjVwcPCC
HwMLK9wHDPA3nTqxLQteac45wnsmpABL+nwAqBtsOWdbTnooWfgX5z07V60iBh4FwUm1Yb9uQhEM
jGhz9bYQuyZob4BeyaXNvIFyfcw5GoelsH05Dd+EjfJxY8zjNmG+tvdUk30MQJgPRY/BNYPliu2s
sLljaZSHcIJ778E7CVZIVvllFfw+tBkU7sSVK/itkXuWQSc7FVSG9dLmh+EbROaG7idmXK2x09eB
gsDZTFNElPBn1VXsNgnUJK4vySyXqAnj3jIyQK+QRaW8sKc8+AnTAnHWBwwXyXU/MK8xLIR6qW8Q
7VvZEVsORIFj6WmuD9eLLI9kiUwGi/rIrQoMO93VbSrAU/JALnyRQvbpTUVadxzzhCjTIXhGsKGn
thPiaCj1vGxp0A3HOX/fz7soDsvhNIpxFj2tSBlbRu4ZuuZmdQ+PbWL5xmq8SRf/lH8YTLwLny1N
7D7FBmByayF8ahdiJeI7K8ogFhC04pVnWbxfy5du/uQ1VVYTYCMv+M9G5pew9phH/2OzdekkbUMh
NKmSqx4wCbuMkT1vUyCFW955MMmXsut3+mDpHpHvRf1jWp67uUYZzOKezYJlrhDae51HnpFo5WWU
pqd7yh5d5WyomQa/pFygQUpiRctnNHLTnXS1I9bvpW8J5ac6gR9kVKS3FP8X1TWLzR4ALk7hrKUC
bJDj1N4nBJD9LMUX7litovn6YY2vR3Au9OG3GmoUw0hF6lAhhtLQQhjmP2QdmZm/j3Pf9LHNxWli
rVNQZxxebko45PJqrhxTt4NwqJziyIfMcR3EQOG44lDhFyTpU7SaE3y7j11396YU4VdaENkC8x0P
JAe9RUZSpcsxE129X+RY+4pFLWdFS/97mkpwGBfaRPE3CsEqzrrCTGgqiIb1Htx8xNqrG7mKDwwP
/TFt/IlXAILsolB9ONOXgjaHgQhBUaBQKO5IPO2ZiYvV8upR5cQq0gVWjmySj/rQMiAG3JTkmvov
1JDlJ+oB3Gs8gfHzOVN4t6W6rQsVfWqof7b6ErHDCNJuTm3UAPBs2S0/uZuMXt0+V/nrbutlYiGL
RBJ3eW5oWYJp+M6pauubOhIE/jzddaObYg4yzRTJEnSlFodgrfyRML2BL88Hx0rfEsuxxuJ2F1cV
O7pzzMNRgf2xGSSpVtOstlFAHXHhpvXiczIl96wXhr7Kf+n/NCGda/nNi2jjG7oFfnHTwc+4mCUP
ixnRxZmpukei9RAFY//aQqu7QMhVnmz7C3UPQaiL3oAS3sovqNbkw4uIJWtCR4+D9yltO6UlmONN
E9WMseTcJQlY0PHEnxCkWxhFbvd0bHM3bxa9n21sjpUlrFjR6M0Is/qYQrw3tVHb4kZb6dubViiB
AOIEPwciS4bMxl82fHZsbxXVGpsoZfRc741eBoUNchcaWQ38PxW5Qr4OhclRUhox5qFTFpyFRO06
0tFrqfrRrpcfan7o1Tpa6hqYeYWsBmBN7lmdsQBaiLT+m2ZKYdH5rXUF9/oRf64FI97IyQ9RGjaS
NZ8wbPYc6jxoPR816ULsT9MBOWTQ/hZGcLVrBi/N4qzFJ2xQEQXv9BO5ybQ9c5Lkyf+Qr8L9GvfW
TUD1eYhWjXoSBE+BIm1VBd6uOWvRV6fSGWr5JwTtLzKjScBjSVJgY02aOn3OPHQP+w1Z4iWWDhIo
g3jmZKtOasKxRi5sry5Tcw6ZMZGtu4297xdYumL3q6onWDh1+P19QGAsT9rvzkRzEWz70ENt0lvp
s9B9zgJk8rA5+as5iLpDKZ9IHVQFKoFwo8WseRU1Fxc6LeLLmqqVVV5KszYLGEvls5ZDLviyaBx4
kX1GpYmM0Tlu4AB0n6Y5+HIdjXAyqbOFpWATIW9CJsmzVJMUNvnTiJGNrbYLIYHaORZZpHp/xKk9
QsVlMq6vZ108FBxJw/8bjHzn9KABsOSRDBnxAwY0i+whkWIxfX49gxyRgy+PtOg0BMIj2lN3BlG2
m0IZ+xfC6Vnq8qNZs4F+BSLNd8LL1y9PuDq0Q6Ldr5lFki6C0Xbs/gX75V1D4AwJOSJ83og/iVnM
TZyKwjLkrHs3OuIvxn+GV+yFyLI2scIfKre03Ok1dPq/brdWkIOjTqihKzHmjB8bYCvnX3ijKvQ6
1l0H4R2yulS5P38ymhbKvkYyZi3rY45EHpLmjA3Q66a6Aq9Uo1MKCZkL4sfIpgGoU6N89AJjKjS5
z6V7hUrsxKGfpReNbCTCTBgW3Gu41PeaQIJi8lqwnGQVUkiPFcU41he5O5+Vsnv670HOooeaF4Ey
Ce2BmbEoo8Sd/MSk+0cFowKI8B0wPUcRrufvR4ollAcDEzK3qKozveaIVDYDhABahiRUUr/ZHz5G
K0pwUkFyFlxkcK+nLbEloY6JzIe9xmqdlxDOMp6qqBmhrFPBgzStH1gOwjl/F106WsOMPTPZb9NQ
AnE5SMRBbsxgK56kcQ+fx09JfMMxVTpBuYo/Xx3BlWrqaThZwZUL2a0L7SvN5RKBAqdycV8XYPgK
jI2sZyomoQGretbsjkTVfkGjoUdRo09wVMbvGnNTMaEJDjRXnaomu8Jp24++2yA/a7rvaXh9GUBu
a4bMuaOx3CR40dpkJiMONe2+sLxasNBaZDn3PpJBEMRKv+tygkR1NO8kcOiIvb7TiQHXljpwWF6b
6WOdv2BQWTHTXe5IKQssdzOt3u/zFSkbADKo7N1rMqdYVMCHrGNzM1rZeMMVyMQEA41QprjJ9EMB
vOwmc/+rXPErjHTOzw8WSElewdTeLebiqP6ZuxQqsA8mHFvxAW+4Co3rJoYSv/W30DChBJvhZ7qE
pvdgLQLZ8ERfXs3gtpgKX6teMucA256XjKGGmxQfkDk7AzmFjwBBGs0vbhy+RlFVbK/H4Es1GXeA
t439CqKnjPSqBkbtpha1CHKnB/vMjHjzgkiSKa7tKokLQ7GCg/oBHlfZ28jmkkPPZGbds2eGj/dq
mXFEF/5fLbHfASTQ0RaN3UhrTq4NcENo/bO6Jch3ec51NHnavrCBvFhN+V0P6wxCFbgZRxcGoJ7X
OeAqqf9Us5aukL3Z9utthqAvz2QKMo+QPlskT5VB0O1738QRjBfKeMMud6UtDt0JW0EHuDD9T3ML
5INXd/3fX5dukCsO7rBowUSvwcj+EmvziES4wRm9NYRQ3YbFU6bw8oEQKRx5ESyZuvDqRItP4bXW
P2iZmc3dIdZbTZTO7jFxciho7k12WUvxG8G6kzbFsifgTrzuw0lhVKGaiw6u9IFnFDIj/ZfVEAjE
hcvq6xKvW/jGLqGFC/Qs581WuCauGa7UFQJ1E0RrkaiBP/MYbvoiW2wK4UcfmSLv1Xwlo0ibQpE6
7wtgtVjT79pQTIm91740rbVf9Af/CIDP9nc+QjqiRV3e0zmWq+i8vt+a6W6NEcvI5cMU0YijAeUG
Zcxbf/+Rc5/wMPdpF7Bamjovq8x23kr+73CUv35zHD3IUe/q4eYBe+NaoJ8Ifm0ERQyQJEsF/41E
lym7OVUjb9ESEtBhGf3H3aeNWoUxN/cC1RRJzkhhBLhByb66iJ/2tuuPKeimYQSbyubsn0cYfEFd
rDI3ZlMX0HDvVQsy/dkkvdXlNtt1JS5NzP3WyK3z8nmXW2RVEuLP+P4/NemyFyedPKU1BDBHlV8k
1GurF7CHug1STvz0jIMmtgv6Gq0ZGV1tCCGYv1HoDdCCi91zsAo3xAsh4qsuLQ6AFNgmyEt+5b4P
F1CC8YkJShRl3Gwd62JzOwkW/CqBLfq/uJTqrnh9jvcTgPaTcpYAtGq9z9Xc3EpliWpVcK+pBdzm
9QjqV7zmfIRIUVh+v2GALRGSY30QdAtGaQkJP07mqB+AI1RZj9iL2M/s7w19xdNRPAZp4QbsAbFF
ZtCVHsXG8Zyd30JHmDVa0NKKmD84tcjnahgIsi/9Pp1ovrSxRVws74kgdCuZcytLzPVsErFD6LxU
WfjTrrRqlCx2RNLd+H5s7uKpIxPK8shzc7p0KsxSyPEzQ3UHH5J6HkqHEDAFkSuJa8AEjYA5ZeR4
8Jshzt3aUJqMyVMgXwcx4Fjza+XAC8qrOTkwkgGeWOe6TkCSh7JidjTrCzZWgXP6qqr70P3avmMe
GW/fqxiJN+eBAqMEslXLwhHjFo1q0VEzhoKqLWp78SLz7zw+doJPVpxREcZO4jLQVULlgmQrHI/v
OHxUe4fc4wNyHU+PW3M7+N/LnWEh2v08yv3Z0vl8TJu2Yj9mtwDgh4bosw9djoQNmPIsVZmHuQG2
auuFuctpPfZoEDNOajsvpDLtY1MtsVZP9lQ5pGeb2VVs7znyJ6MpTgV1HjSTL9ESdranT27maV+r
3Vb0Q2UN5Y9DrncOgT0WOyD479DMvkAqJnNkOeFqc/q/6ziZfSRKiYRRkCaNA8izMtELkL4/ITBX
j+I55OrpnDg2d9mxWIyyBv1maEWMmEbeHvVf6PKIAEaHIuMUonA2RagHkUxWY470wIbdzoE44uyr
IsZREbJsCd80DoHBEMv72ldvWuejJKbwQ7maW309aomUdFprfwzrjDHkQgMNj6sNPp0HDlEv6HYr
UvwekbiPXpHretccaciMvPQmqlH4qXO8xiTy4qPC2DQT+r5k3Ld4W7CObrU/UEarfMCDjW6D6rVU
sfZGMuElrtAILFIBQUxQRF9qL+qjYjka1MrlX6Cx2D5KVcY1A7I1O4L7Y0mf4qfedyogzuMUNL8s
yqFEzbMUsXqEhV0GO+DQPyRkYPsLsKow+L8dRG+I08sXjjAdycuilcS5IjjUHeFOiBepgWFA0+Qq
nvc7NIkeGBDNoDoxQeQhJ1qgDMKEda76kvE0z9Vz2r0xTaqpR1LPIu9mBO2hcc2OhJLDBeNhj2CY
aqH1ddXkiB2cihDRRxFxfTyYcmOigitrSRfd1/T5tkay0AKPydzZp7ozyi/Pz4tTureUWOL+ap+R
a1vF3NUcx6yVVJN1qgfGQ17dMf/2meM0AetX/shJIPtxJOVh2YF43rUlT3sUxsjFZ28wOaUVf243
b2AKRwe/i3vSKoCvi+g2tRqWF7p040cgQBoRqTtVFw0yoh2WUzdeU4sX55B3w1ZuFuLTr7WWC1qZ
LlzlpcoOqr4+VlUoM/Evxm/G666abrn5/OjssU0urwV5N12nIqpS8ieqz7WZTj/U5UZiI6Q8fMTD
vXXSCR2DUwxCEgysuRGkcxoQ8KBjWLA6vJQhr/Ck68Y7LMpfiEx40NMt6nFaCGoyGhQ7O1aZWhOZ
NyP86FSYudM8iF9YOP+NrgtT/aiiPjdSfHyRumHB6ON+iOAPOI7ulEWJpkmPEnSETMVbli44K95l
CfzppRy1cASf7SdTUgwbhx26Tjw4kdBhvTSVoDcrfiyjOMaraArD+CqmMpo6Zq3XwK2Rsmon1sZu
5CzIZiyjAvQio5CNTmH4UowvKF+EDkfG//erpENq7i5ak69UHn9ToBETf7dY63SEqdtc1gEQGz8f
z+NLsDmBIqvOraxX+ZXJxjLF87pl/K/kqr9NVWuu+ekmQClGUKe8m0QBQKtPUmI4LaGqf342BBZ+
2gFJCP8r8NaM6iNDJ57UmHmBmZ9tmbFRFD6dUR1+vOppNWlU9zTFrE+QocFh5Z1SYpiQ9V7O/m7V
AvHNaCD9gE7BTKvJAvkUdWOD5KvtvxEwI0w1G97PFQZC6FbLd/TQ51WVENqyd+gTsXPjIDXP+9nM
3m2ALA0ZyLKZfXCxx3i/Lyg/Yzd38wd8RlZvkhLzFLk17GnEtMz8bueazmd27s27YgXJgTs7VdB+
Mp/NO4tjecEf1DIwLtup7WHdZe0BcuSgMnu/ZeRVOwu82VgHNfbiNXC1pdsKNcTg5C3f4PJovUSt
iOT7CW8ozaYX3I1R9qU5w5/iaY9j777Fdqebj5jyNdObwszsBGFroaEnAOLwzfSGVF5nGa82Y71N
LPfuFAKB9SnzaJOle53uP62aNMAr5s64ZQ5XXClaDfGAxU+rkKjIAodKp4Py72QGlmMUKgxo/3M8
jaYFLObzk1ZvpG0sXgfbxv6HLBucZIA7SI6QpWVXmAjniHWe0KV7JCdAnmtu/SISB8WjmzxkfmWR
zba/AczICmBVPVzQXGMLvaRW2iRJ2revLYBLZakbEZSq0SNpOj0DfCloKL4ev7ZzFkSCUFMa5Nr+
DYESznVnFRGbpjVZwSctkZwcGXDfg7jV2I4yN7d3P2eCVJqAGD4rsr+5KizPYYltWNjcB4j1IBLe
YFadJS5pw1tpqKym9Bn+DyfjTzo/Eg3szYLh38FuQWv1hjBM6SfbQsI4OlmD9t3z+xNc3N44uwQI
wswLKXeeoBGqFYzDajej/0u/NOlPWhC/HiJcPiX/WMD/XiPHTQRYYMXcx7pSpHbsyR+YB8/vBG8d
mkVh1cLo0JDX80UPPFsLVEEq23+kzy38Et0TK9bgMBCC3GDWRAve5vMnck5EHW4NZTPWnrXw4l4Y
iKgxy5nB74U9v5xL+HGdd/gp9JZpFB2KrwFl5Ng0FEL3tXSf4zlbkKFekejldCCKREjr/D7CMN/J
onIUb4IM+bQYrHfetDBg1YJnsXdtMgjpqxHf1ila/IpNRKS9aegGUW/wyXUXcRpA8WxgKwpTTr3z
piUZ0i5ukJAJ4t2EXjuZ6xzDFHkzx+1t0tXsQNne7XJhFAzUHnhyq/wfPs57qIs04BnTi0Qha85H
STf1vJrcNY69pkMPly4xpozjGQ1AM0gGohADoD3Mymm+eCe7ElIXzSdYH97YOPz/TfQSPRgRJYa5
AkNgSV2kLJ0ezZWjJjxp/O49AnUbqoEbxRSa2fk2vOLm0xWhkIxcSozufuitzn4kk/ClP5uxIDjX
YI6ncHX/c8HePwInLybayrrvskzHKwAN/4uyw17ZBejEpoafNeOSmWFXWj80yii3HdXI+asmU4IA
2IebY52hGOYkKdr0fu4Wu0IL2cNa0/WMtsVNCYAmWVK935AbX6Y7oSKbrrvespyMMpxne+H1CKrb
lyqev+I6uArC56IpBa1KE5UaRANHg3Oke/BRKk39tEpvB/qar3KK5mbsx0tE7EbeSlWUxByPRmku
KGZ4mQRuxPaHT5+lTcv0cjQOF5uiJ37gR0fqpSQJyxWaRNjjbbHpxyxVJqMclHIC3v18L6E9tkSj
pxeoZRYO+hzOl7D6rnzUyqv66cuF0cTaD8W54AInDkLqpSTjRFESJrbMgkZS1q+efs97ebXc5ILG
XDaVK/TqmgcVdi9pDd3ejgbLjbqddfJpGD43Pz0GGh4d5tVk85rke/sGh+b3v/nn8hTr9YT7QkRu
Q/DqgPZsX0lUZhR1wumipvstCwgUk16v/2HTzA3+bZM/6KrhYj3d0vlnmUTPBV4rqvjhhxvQSJZb
Zs1NliqCGmzNzU6g6dqnVOU4frNNezyMNWuLnNtVr5W7GQN9XQvOJPXJDlbZ4X4qUl0r9QCg+UdX
kFIvajBTt7CGvv/9GS0fNCPWIncCAMyl1Zk0mqNq0YBZAsn1lS6LoIHNKsQYQuv99RYIDzx/lpXm
whnSmcuLBuJXBWfPSYgeRrphcHHLw8lTGt+OHI/FtJGbjDMMy+6R89Y6qMfub0cHs8HrrYLM9jql
Jk6x3AvC3RXuFAV9WRPYa4tV1Gkk91+Ul4s9KRO4TRA16paDMGuOJDs9zjhfTOlGzlxMUrBYZpjx
Q7KjeNn9lA+YNZyx7G1x3eFCRSWDdRtfJAVAaXKRwGs9KZ2sXHdAGILFbp9akh/IFSucTGwu2j45
5PKD+B051Oihz8+5hePqQ9iXIE5pAYCMBqNur1f0w7IaENKfKuTjSmtXd7XNulJZVAU/U09aU94w
GUR5dcY17QgL2cLkr6Dr5nxdIngzkqCXoXyvU36K6jq4l+/2OffL8BghS3JxJcffarfkL6WVhhhn
avUKDwj6KDY+W5qO57Hwp1Zg5xF40iG2RlEz37XdqIt1+YfPO5mxuT/+P2Bhj7CUrvp/bhHfAEDp
VqL2Zi/o9IHN2nXUuuCMV3jvpvNMZzNnqI61t/M1hp/jJ0MkgxFgEn+XWv6MHgOa46nxMF+zc4Z1
TMGnUx3AWKi46NlRjirKvQxO0StgxgawkNjo5qS3Fe7xhX9DVPWYjnIswNnSqDN5/9brD70zNQKG
AOOiBWzqBt2ROZdWoUGtkQms3ftNYacFqLE5hTX1lonD1Ijuqc49JfK1ZKrP2Gqf43hhwa5R5OJY
0iQYcYgLRIRZpDV7b3fpDWARHN5hwoilhK1HHi6XkF+upycB9tO4cQ6dX9DauJ1WRhvfvGxA29Ji
LGV5fI9kzNcRT2CZlB0hn3KLbgORjhVqi75oAOIo3wrNNoqHG95VQTiObUXCw7LVS3rFpQLzmT4I
nweXQtJLlfxnmt0AxMhF+E93kilNcacLpSkt9T7IwiKbafvg5fuDr3H2V3TGyew0Z64q+AB7bqvX
MoLY0Nm5umviAI6iFzF/2oM94/VFhNB9ZG6yoTpWj4yl18/tTiA5Wtof3uKRzBj0u7xdGMBvD47u
57ojUNMfneKnvs/weNgrPbU/EupAgfVXtGVoKKhSr2DUbYqQ8D1twwDsY2wCTaDyHugZbwbHnpwp
iXJC3A/cernlahFl9Sy4VYi3cu/PzpazPGJei+EDJ3q8UmlS8MXG0PCcqDNEGVz+JO+WYX8c6hWu
dy/Svxuhze/juXeQG1TADqVSRiddTzFUPS7ezZM1H3FxYNGL0OYrQftlQYcvDp0qSdcXmXV2K3W0
tqRTux7vNYhba9wHoqZ29yptjDxohjv6Df0P/lv3U+cIDB7OyGfaSnqLDlyFMhkCOmvw6ynnRM/t
q5zChtgtyS+C+vug60v+/WfHYMv+yPapBE2CTi4qwmxhObc5J5KpZe5GTHcvVAYnsvWI7omCdSy2
gZglf88/TXtLHs3MGBKLCxedKB3HDhzPAVQUPgSI0gg5EAivdIgo1l+95AusmWgJNkVpHPd2lbJD
fw+SfuOks7+3Oz1fLabxGAE8wvO/SUhlGCIUqApcAWr/nYQxkKXvAjyCVlLTfnNPxt3q1FayqDU4
E5hhtA8E8ededEf5KwM34J0YINufBEmaGvZmnNeBvz9pFPisNMdMzc9SyRpWQtb6ZI2zYjMVXOHX
mp18Cm1BkcfUfab5viGH1VWadGGpXzwW2VMvOePnqFFWGxkFbw0NCOtiYKwbAPU0usZ3V5gaGXqi
npYBjbGoZxZkffP6a5e8F3q2aO+3yfPeImMChDCJvIfCNgYVA6CKj48S8SecSDItLkJ2vIOsF/7n
E/XH3QD/LSgaKxOetNBWTJOLKMLjnQ/8rL1d/8x4DDKKURbbXkquJfjWNuo+6TE6HZxv4n28+iWO
W3dk5W4nT3op5LEdXi2nZKupdxm6uXlM1G/iJT9+2FoQz0lI5uKcxjTchDd/9BnJzks7BqzQqBfX
BZHXDLMhZgBJxxGkCNulUq3lmlghc6Nr+/hxawevhK4p8ArxlETx7wUzIKsM0J5yP/L/0y0VQLrK
eePFlo1eVEsAnz0giceEZSu3UFVOudL9bMjrj6lHkAt93I4B77VYJ/dY6CbyHsFk8VUJ4X+mMe75
psr2jc8MITXRLefOL6hBssmXOFV88in5pdS89dq1xPzCajvK14JYMiUTLggjK00Dfs6piRbx5R56
6AMr2TycqCEIeTvjO+TVMmig3EIKJ6CancMl8w8DJZ2G2kmLSk2NtuxLBtM9w6WyzdSC0fLQJ8fo
oqkWp1ln1muzseQHD+pZGn5eEeFoaNvg054kqw25lJVrsTKX3PoHzLMVPIv34pHTzvhOatjhwc1u
YiaqwzJk+GUiGDXi7qwFKl9ApSQRdrGhqc12pb5M/Rwdb6FCtByIuGnGdgf2yW5BsBQdfLrU2pXg
lJcKjYOIa1g9qvCdicMqn6I8AjqnHMc2jBfsHIgRONyh+cRlCZvdvvpZlxF/88gfqS5Vw0Yrm6ZM
5r1ymWoaNn4NlIyHyiM8pFd9u15P2YeooZTB+cBERB5B1aLKnw++xBX+2kI48ieSwmDN1rKKH/T3
Uz60u62VxsQ6xKAYF9zWLP/kVOCFkJi57jO70D5/Xw3HOTtxkR1pcSTCHfwLT8fIXGQPcPRA2ksP
2fesbk4BguxfhNfNMt94O4pbJUqOjQ6U/dqvC6yRqASd8OUOrLn2PkRi7VEHMq35eEYbf+WK+Srt
F121rroXYi7APOZOcncyMRNjDQAYfbBHvpspjxO918XAysiIfnvE1aezk4Gpze53iov9aWVtV/nS
EngymrgMZKwBnRB+cfdEaIMEfRdzWEzqX68B5M5f/EBrlzdps2e5rncsc6vtXaVnrZxI8XwFeXqH
KCwdelaJeNOxjKT1lrAOPJYjDg1zN3djz/eUD1oRP6xxyxoBeJ94qEOVpUOTEdQz7alr8/xTs+oi
yQSD+mq7X/T398mZPvAVtXq1vwzabJ/uybOuD6sg4UAyDHQOsRePjtk1PwkWzA6VXUHN7eRrUc0v
MOEl1AJyuC61bs6e4ot9pgtOvEzM5qObwwCFI/l3b/NBbSKMuGeBZ39NXKMYmbpBWmaebSqLQh2V
XADBBolEgUBbm5AtBeXY+gY+bzSjC2g6T77joIR/8Mv8PbW6qZ1vTyBWTuvIE404yhgqbVDpehyp
7iJpqxDMizh0xISsZCZlzmJT11jlEJDQZ5/Vo/YpiPl8UKGoX5MPGNHe7fnPd/GspnW7TUXxvkjJ
tBh/yHkIrcbwj6eSoXe2IXI5xSMvFQyYU9FN0s832dYDQOL2ESdT4J4DmKpqjbf91U8JuK/GwXl3
ozNm7nlze0FvQSN8Hc0SBgot1p5ITnhBMOdPcU3PdUkcuofmh0XFrjHcw5IGTwigtVnxWpGs7sL4
tgJkznL8NatKM8ba9ahS0efESE3QWzK4iuh/tGDjp025uRZIRwZ4GW3LQLv9UYdeLK0epl7zUQ29
56o1T+ip+vL3mWV2ez8ywHoZyULbM0KD4VnS10+4AI/ckpq+qG5wy/qy7kIRVgDzIVVn8Cls80IT
J2X5T0N7bDtcJDpS8MH3Sy3nX3UkUeqeVziZK+hFPomgyDd6tzHg41HxLI8YGpG5JVK9QcBLvYmZ
9RxRFcKLARm34fosLePlI6Aqdv13SIaWI8VauGBJivhIHJuRl0WaqkrCau5ho3YFYM8MF72zcHQf
ViedlyKKHmD0tJuzI7yi2xZtRcFZgOxjvDWmEZOdR+zDfx3gort4Q0tEmSMAnRXPag6wRU2eJWpU
OFtVuzWYqXcf82T4uvPIJ8RGqyweKvy2L/gixy2/Ql0XHqgwRhFzyInF338rxo/QgPdhxOAByfew
xF+X0xpZ9vgva6uFHwUl/UmyukISdM22ybwxHqxMvDMKGppvGBRUjuQedjQQoHdJS7QmqngQYJGB
2xQXMlw2tsqCN6cpHtZwzAGQURWRkr+8Z8HnzhpHSVNGbvwPGIn7bJfpsu/9u9R33xkSH+ugR+Ln
ATyucSj++tadd04CRM+n2zi2RuRMWZ9qLcCD3PckH1Tchi7HNWirNZfqBwpQ/aL2prO3+EUddtUc
/fzqRIZDUOybNvQT+n8faiJ8VsMtgrx3kxwbuGMF5X5wbOUUQwBzAjiygqejhBHNsk0MshLhpx4T
eshqZaO8kBC/wx0mJbGamCKnsUfzemBvqwLJ8ZfM2IPYzKy/FXInfe9OERt5eURpV/iTmoJfuWne
/4ZnHtLGl0FWRMIiWlasAk/KnpE9VXqDcT5PGcigTCC5Dt3lBapgQ3BVd/YbeNV9b/enf9ET7raG
uHyQbvKlvDZl7ZJ6zLBxqrdkWmZKbV7NxDqc1urDaEigtVxtSWGorN3PDd7eR8iDUgQ/FRs1cqHz
M8gKedgvscBjM20/gSxZYfDICWz8RVB64zH1YtlKgz05Fb1YL2uPETmqSKJW15Q53B+EDXxcyuA3
iQ9qX37gVNw3EBEBXn/mOMzfqtRVaQxnU8HIOum0DD8YrHEMYZ6qsYRRHhU6hkJvJM/q6KNiREgq
hMOgxc8LYvrb/b+Alz6o6UPl8c2sEnf6ddm0VqfNs0AJKomcWFtm98ERKkcWhDWh/Lh78oxuMUpV
yQVu3v+iWGO/sO1yLCuW9PIUqoYd426/1yNTV8GLXPsxO7U9T++3csilQsfOCidwvpLWpAGu68cj
bej6qAmik5F6GSLWn/5+g59u93wpXtEZn1070r/H/dAa/jOjFv1zJ5fbxEAMVDDTjtz8HbXRfWI7
O4PMP1maNJCTVAoe8/pNoWOKS/eNKNpq+QCmHUSrgKVL9qKakGRQJ0Dn/U1WOp17DmWJrOiEQDuL
TCbaa0Xla+KtDI4Q7eb7CadXoCH3L+06Miew1PECqW+MUIgHG++eohWEPkxKndVc2NL8eLlyIuJ4
mZst/Om7WVj0eB6P+YzbithSn6Sl8paUFbwYOQdOHwED17jwIJHtSG6RV+PFRJM4mBCkk/O+bzsT
xAVD/vt1vKKLotO2AKJjA0ZqA7LUWwbsVQFQL8cSwIJB0r2QDP4XWVuFN6G+LGxC1KkNZ596eGn5
m+vmNBmluTTI4DfSaGanh5Dd94TAp+nKBQ3CbIWFLq8QQ0nPN9gqj8CeXUOKZGJTFAu64N1BCbeo
GsLb/OyhlPaXJ14d/zW5DEcV3HZ1+g8i/GrICvKJ9cFaPyBxah9PElU+HInjzkHxoy5Bmoem1aAB
EZNsU3FId5OKaiaL/TWfYR7o4okw2KngG89CFVsP66iZnhFB3AT6+uRZKx9eUH3GQnAlzQpMU3vG
SzydqN7PvTQ0i7IA80BGIY6NjJeJ67IET4PEzlVHpbXjJ08MKdq7xt7KY/IVLZP256i9s1uPJ0Le
c5ENIeSS0S26bJS6LOi03EdezAzxpwHiGj0rbIpFHXoLK+mhgjIMiEM18aZm1sCJM5QAcw3NRfI0
GSUxilV/WuszCjUjKRjkJs6am0a9VL/dV6kZuQwnR8D7tHo655J/t1DswWK4CXmjy+N9PDLBdg0z
opQiQG+Th3jn7HOi9ABGDWJATrsyMhlDsQrOLfwsv08M9h2X2+bBu7zYVAFLpLDZlCytJ1o2tj84
Du6A8uvwcUgYzpMGMQ963HuM0EJcGASqci/nTnPp7/uUPxyfQzEpU7HLsd88qkzDqhCd92mJga6b
k/Qa8suXFNhduB8W4YcZNIoqUjRzFj9ikyc78B8o+H9JuyJ8+zRS8xQZiUcI/uPTYtoZ3Yt660MF
NSYi5hyIdgyIOpnhbDMO/487G+OooPkNfLRrPx3Gzhan+jPvrM4oMQ8mBDyIuUG9uXGmhvNtF6/C
GuMzK0tx8J48TVxSZw8bgCc9+1mV44k/U+9SFY4cqNkNPdej1bzEluhL763zP/Rpmi9Vv2uaFe4f
OBIQA93wtdGTDoINjSp8+/ZhErW2SMxI8SVSWOIrvkD8i80Ua6awzhMB10aRqYRwM8o8dq2+IHcp
x/NFXxmO2Xe560VnQ6RjRH46Xp1zXmWTN66/ztl6GtG0I1zeGFYt3yCSzlylQ1QBY5Tk5QKcayos
cd1EPnIgOl0Bag5yvABJplSuwPNSXUq4CaR+v0CCBmmjGV+LYe4aTMjDO80l7Mtkti9LQz7gU5RN
kGnHYkl7OQx35uyhZe0chATRX5tzJPxabpjn+Eoksn4Qr0/Xh+xORNX1h5l6Xj52QwlOMzUs6syX
6yf/lsJoXwkIjyOY/vlZZZvX18sfITH6gpTKpBeenZNz8UtFu6/2KKq3KVU704T+gN6XH21HzQXx
03PPiWTrf48KViBh6txcsIqfl9y8szFDHRzS314hBecLDQ5jtO3WSA0S0MpSYIwmgZ8TJmJef8K3
En529BMYpQq6VhIm7ZI4QudBejS5qmRLHx2qu3hfgXzglXLcm5cXmmgQmPfv07UZ+OxJ8xdbz+rH
pZU+sKK7mO7NL7pXrIbJ2jFy/LUiKk0J9PmeumhSR5gRshf+7/0rNNzctETi+Zy4ndQI1sZkR7vX
DldyebHcdaJ8iTB6/y9bkMp0w4bzaev21AGN9cN2fKDNp2gLsRSg1GnqTLDpAxUrpsaFPBzTJ8P6
grzbUxFozXaOsRY1tAD08q1sY6eS3DKqbknM0rGRg1frw71PPcGxyoqoSqa3YtWzXuLtWbN3aczs
CteX/APWdaTp/kNcmf0dYDTEEaz/vyugFZvPiqVca8GuatVjjRqYVHBFu+XwK6u+iAeHtVMxwLMj
ThhrRGpoii1zXmAs8Li9UWkp0dORKvc9zTqON3Tlmn7oyu2+lLtpoHfQsFI0mUT4NgaVZHY52YVg
wDp/n2VYBSb/ZIE8O+R5qBmx7HSLA8TaagTQ6UEtK+loP1ygmPWSqG0/OwCsWpGO4QZ00wEsBSy7
3uMNvjCK5HCOVUD0lmcGHZGvvz7oF48y3qOGQ9wHhgEwwbdgWmcKNWng9SO5j8ZtUjJt3SRtHDYX
X0ll5sQCudgSzeDE21A9i8IaspUtRrRa8VA7ScDsmO2fAEgSqtkSZMchhotufaZASS9eWpPfVUMK
Zdh1xS7syDdsdUia+7OVhXHc397eWqwLOBUwfzOYsuaQ+NKrdRFjcUsxgv2ie5oqVPdmSUgGf8Aw
KdPyPNaenlrH4y/o6q9kgMeZGZMSF7i8BQV8cg42A+FVHvJ6WpQcqQBaEwKugaHuaMPDH3JqdXJB
SxpDbprTddlhR5dUOMnzo4L4aPEsssoKdd9rgwz/v5R59Vg/MH0P4Sp7+rmPZhHTbkypx2T+rv/c
bZmckw4jwoQjHMUoS46z3/Ho0YWe6XQhKjnB1OtaQNMTDwPxNqVRrPBq1MWoHIB2z14p5UoMUpaB
PLepKf3DwWbH6rRiEow5jXH8kmP30KY2QUZw+BhOo+p3VgSAtMZc9FKg3ywPbclhzk96kYebuyWx
mB2BpmyuEACljZH/foDkQRRkLXutbqLDXJREjrBNxED0NbKPeOi4asok3GH+odw7Z3aQkDXoyPUe
Aw1Fhp5dy0/iDQoj3Vvpvc2rE7zF43QPt9MX4EqNvV5aNER53Px+WtV/pDFD9PJtxqv2nR19TM5H
uhTXQLKBL92aHOsWyYH1u3OsXY98/65sGG3q+MfKaeKd565ijUuu4vgmX/IscCJwSxzRzf8hy7Dw
aKblAwIVQAplAisb4sfMzB10DT+iwNqqhoQzU1BBoyu6+K2bX5w3hnbaM49pmVh8dEKTDk+lStfh
wJ8z8MOhO4xLdFLklzWOe8N2fLv0GLvF0bHy1SgEPHt3BQ0ZURX6JC0NuLU6YPztx730aDsea1kD
6C8tUhkJoPwvm+cRAx7CIw8DxZ4f/x+zuZ6ZeSiQlMvG7b4tIGRx/VPZSESgzXQdrEKJn7ft3zQR
iY3IBbCBtDIDgYvrALY5jz9D4i1hf/meHza6wLPN1oNeqMEtJVeghRCkir3Ib+EOJiGKhbHSBX8J
7fUbfxbtq6E2zrtdNHgPUlKRRWuV0XBLcq1kDC2VmNiXq3QyeEL1pWnDQRZTjeswoVi2OJ2ofk2a
mA9huKv8WiR1A4ZwxrmpQe8FFTrniJX5eP+YtCHOwJJ9M0QYEVCibac0jPR4ie3WBAK2Vnu9gsdW
F6ebgvi5X79x1skqdi55aaN0W8gsEFyhgDAA5YEO+IIZq4c74wgSByFZzWhq1bhkWg1Ye7c6BogZ
np194YvieFz5I+KuVTVtoGhcISLJYLkH743OmCU7gDTw89QZSxO48AoNDrYuI/gkv9crKrLC49i4
FpinKJyfE7a+PENiKvtRFxwWMWlukwL514R3hFSBANsDYztpA9FjAYEkSOeY9ZSuSSS6397xEcZU
QfXIPHNhzATEPPYh/igs555Mz1ZBt5BOQX9lYnGt2VxpOvhHVIJn8HfJ9nuxe4+8bpxJolSkPyrv
BiHFhtWZnrk6qfyOhLPdDCUSTv7bOeoNUvQsWu93t+CpWNtW7O/H95s1QqEqWJIMq0BHouknv/IG
In8mg5DdqhttCpwjxPR2AjRDVZvWeHnNOkEEKYRlJwlqqbnDl80FFSdWfnt7VvQZV01USFp9EwUo
yOBQUFSagVBKc/uY8wf2D/gWZoTa1lb+3uya/QwnWXXh07EvHWPQk0mHf9Z4HnOzjD6WqgOX9DmQ
zIejYgUbRA88ru3ARP9C7Q/oM08a9q6M7KDCot8HGGuUBxi8o3ABlq39sgHEMKbQmSGQMtkVLHbf
droHUvPBHHljO6Vuiwl8pUThBHpQlBtYea7hDojttHJHDuzgmknYffG3A9q/Q63J0QWvZx3vtKcp
Q7XXNfSIIpY70HAWMk80ZSxSdh79aK6br0u0KS5D/UT+YF2psipp1telRzekQNrD5mUGeCoRKp5f
MLvaGx7uIGnvKoDij1pr4BO/LDncCVCO60bESHs6EtbMO917PwkFDvcDcdGr3InHv9k4hcgtOygd
eWNp6qmAg8qx4Y/3Hn8vGxwfTxUwZoxnfhcOcTN63AHqgJdsKUBx2nHXK/a5uhkOd2n8WXkpnajU
yr3G2jA+8RKl3cF3hLIp5vR9ZzUBJyVbnEdg3yLGA6YlN6lGm1ws99bvJ2sxXKS2a1S7iwV6YHHh
lFDExZlj5rfBNnMXxuCLYVsFWtzwyORM0SjFt63+uVy7MyBgCswSVMsWK9YAVN8r8mb3W285oaCB
c9hFJoibp6v7eKJpKZAkkd0Z0CEae5lkt5bb3tx7mXOKYFWBHEsznHIrkrs1xYrkqh+ItWn0VqVs
zFg8ktraMJkM3cN041d790ZkI7NFFb07daZ34Qg4AyY0NEc7PtKoAnGkYKd9hygzrg+T03MGm+XS
p1hVIcDK82BjblR0y0f+bjaxIlY8jUtMaEDay2VgBHKyMzU/TVZUijTW/HOeE3w6brQo0PqGAtTL
J29BERzCjM1zVintel1mT3fvNIKU2uUMRPZuW9FlFRf66Yg8JcS6+kq+9pRKpvwuQTu1exWpeh8Q
Y15zuSlvU7myHd6mp+0jZualtVZbWg79vcf0Oi/MQZFnX8ihYkqMNd+qfEwzC5d5LIicXhp3KF4e
186Yxaw+C82AQpruuwkyWyX93eFw+GAk/eQaZaxPDh4RG6PquRq5NRLWdBqLOnq6v+CbIYKaKjAI
q/rjOrtdrgh+ueuudPIWIV4u4O7TqJ7e/+SK2e33vs1W2vfDs3M4Cxdf0ijCcWp+LOwSXrn/Pn8C
ptLzdNJnrXID1DaSsvGdaEHHxE91EvgQF3T/L0iOW/gJ49JGlv/3LbwBH6KK6dlGlh29WQtJGcyo
XXTRYFtjIPq8QgI5ZCcWphn98K61CzLiPl/O/UCCnIaRfGmUy0wq5nhvXggNJ8FtmO4Kkw+BN8yw
T7nM8ysfsda16Ah5tzzavgNexej6H+RjssAMRoMEhWsBKf+hSTMpnbrZEUzrJyMavNkM+heoNmYY
zKLjBXPswK2WU3H2ssZy+GTmSRX5iuDVWmkjDtlt3og7FH/1yBMeL7sLKg9xOJEXJRi3wyGTyDBj
ufYSczUfouul1ZPRqmRR7ycGFHDyTOfqdw1TwxZx4GUB0t2NIHhHz3TBrOnah/TXPeAdIqH/zWLV
QRffxEIztb09dJpR8wrxh1zXYuP1BpUceXlnIoGXlPnz0vxg9xxCvAEuoxZFGMrIdCRJpOtdGono
0M0/9NbpAbUCPB6q3ewmkAgaO3VBwp5eakIHSQ/mey0WlBg6JvSHZn3gkkpKZAxJqcwuiIFAmDbT
wWXuq+g8JmnZ+j3XhPMOkVuZZAiU0wxWxyJUKhtimLVY9RhCX+Cn1caKuia1c9ev99BkrycXVafe
jDF6koI9d2m7N5lnj7CMOeTwi/c17HeB3kO9iraBA66uAmDp3zQmk3BASzlYMQVNVM24MT+CMjSS
ldmMLvLAg+3BxS+DGsUbc5d17Ij9MkEdp1B+9552DxSm2lVqjFNmtxPGc4SnUWHqVu4gOA34xVl3
ORXVY6qDg5NkiN+xVPWA+qSuc8px/VcYP1QbDPj5TQy78RBY+sLAbLtX7GmvrsaCInWR4x9c4XkE
mr+OQQV0NJuJfJ4p8+SDrHCfshEz/I7qc+HDATD5tpczKL/B26r5+TbO8cUOvKsOOUd+a4TwvfUL
EcdunxQcPLE599QkEFGi/u2oeOrPYuGAvnoCpJoZslpwhlFSbEiFSmX+v/1RHIEo1zzTlbEoXNCe
utomIFRA2G5GaajDGnPf371I4j5PPb7wv82nkRrTQQzZNAE31TU+RhTct/Zptf7RCl7ZyJAccwWD
J7DIiYMaPoUo682VhPXzXr6N6NjfhHGs4PgoW5+sW8Gu6kghBwOxDFn1K62kOduPP9uYyJXC93Ql
R9WWODZJdDYRmSC8J5xq7W4xGjIXN8NjbWy0MXzbpkFhCw8HT1g2EbVa+m4vUAW1dUv5m51njtdI
GJQ8FFad1buT/t9fxIeOFcmiurIm6g6AmYXO8qa0IHyjqB3BdkkNR49RNfiZmnGGuo1Ri8GFkS7x
A+w2Wq0a6W3oH7FWgfV78lidATmfkT6ozZogwVoQRvh97LDh/bAOh6nMWpzQy+eZ7DWPpTPbf5jB
rcjoR42QQr9qy8VEdSBkCS1ZRZoK+elB4VZ45vJhv/ScvgSx9p4B67sCSnuJPJzD936ZkJt67SJf
AlnTakgXHQVGgjgA1e0Jb+rTHBrIerSANjecX1Hq7XPrmpi7NYWf6xXW3F/NHkU1Frm+oW1VBgjv
5HmfoWUfV4uywCG9RGrSxslATG+ipseXvAV8yjvCPIchCzjKA39cwKyxO2cZrEJ+IESxvmRozQzR
Yr5bcdgCbd9kLhp1PmwIMIT5oG+mTffzjEjJzWGtPWCQ93ixqpBErn9jKptkoiRF+HoBm9AwumNP
1i1wZ/c758xPkbU5VeMWCB9T+gxC5t0j5bPTfSryYvw+c3cBCnqLKi5JPnf6pbrZilSyl574Xh/Z
6vSncD94H/79f3sa3Z1AC2mwbwwfH28g7M35510mQFdwkVY2yXGLj3zgQYFupjcGhObSpkKogIbd
0GZDdA3Zn4upmPCgEJBN/KSERy8awu6bqPL5+T7Nv+4qtz2a0TsARVYtmsrDskNBgeYSUHplBLrs
TuMX21VwPrClx6YViWj3gveNauM5jxhpgwtdnB30t4sGPn+aZGuu4R57UqqK1MEMRb/UIjDT4LMi
/ebvaEz/3iF08vTA9KA6VO6qnODKHLNwDlcPTR2Dvg0rr8222bPKOHQk2NVjvdSxqwwsKeRotY7u
HnsCOTlGx3XPZxK+IgFt26TsGofABpZ6e6W+3hUgt+XOFSH9jGBTNdxwy7H3iDpobzgR3lgwhOhg
WLyNVCGZ/AEEOfOKpkdEWZviIgD1VEtCAbARjjS5a7iTg61IuIldIAxJ7e/PEF90WdYUhbMYrJI5
PnuRdvQT2dWecRbP7gPq2wTLN58qbd+TM2cpXDDPnBuThAEMMdAFQ6RxPPsYbTsweo/zhd5XbWX1
cjVJjOT8u2SWmO9NSu7SeAYsCi/DGpNNfj2wUDvBJJdNbwajqYKbBAp0sqork6L3yb/oT9CCwiz7
DmqyAPXRmL5RH7rqZqmZrL1MVKE/1NE0Uq1gbcUamwzp6H2dFqNoZmWC4R7HK3/g18SphnDVB1cF
vXC04v1+wv0EmnBnxlInzvJeJr/yXjN4HXWbbcrgANvnEdUibtatXM+2VAp1fLBFRsRrq+kF+Vfj
K5eNfg/tA/fyLticPK0y5ZeNOvUaDeFm6U6QuyTLdraOBbIiv0hGBI2GH4QuH+Pofr0tBXo8eWMd
AxUWcf8UzMzYaShTt37Lr5VefrYbGGV7+yUvkYyvJ0GoBhKeyXubMokKj01xJ9pymazB4JwmV0+M
86syKk/mv2C1LgCM3Hqp8pcTc1fulOaX1W5ESKR2WfEJMPB/z6ZEATjAgCSJkNAjGB3faME2TGYg
v4vextlkTYwu7cTWKwau12u8nxBP4tG0Yxu3OwoHX2JJfy1ME+AP0OUobGLY1WSDst6kgreLkEtw
brAp8eF/hjkw5PIAEzH1yfETJjzfzRgR+ypKWzrMsltzmd7WLhQ98UxGUg/G/SOTqdiTGjik88+Q
UlimZtfH3Ufttu7x9+lKfH1FBMF1aH3021B30KbdF3apgeF/buiBWQTZzR0ny7SGQ577YuCmICf2
JI135CcOmidmDl8FFLkeKiTjk+1Tn8HTKAJpRxiS6CpDzHH1/ZNHLldbFDmIdfrRMDZFsFvhtzT6
vfuWNZUpdC6VKvp7hz9jTDA88ZQl+wjZXIUF+7b8DB05/217gHsQr9qAQVIRKwtv28O+MeZT3eg2
Pc0pmUjCVvyWUxfiUWoEcwKoXy63c1ykGxWUPr02ZMpydCvGXN6q+l66og1uuUFE3CVHoNxsGaiq
uM7Ix69AfCtqRqk/trsGFt2ugqdLwxty8EGuY8F39x7P+UMttcEDoaFBFOyQfE2LWSjTZGC0BoAD
HdOGSrt0y/2jhaCqEPz2jwECa7Z4RbCGC4e1ylA9bZYTh+UGvNShgg6opBb/8qb4LComcN6R7rMN
1bdrOfGu5pqKc7bVlahJ09V3ipByUSfIhY7dOihiSkuFXynflOPyKRkj3gv7TIWS4nHaChEvd1N6
+/VGroxdJUe/wPYk1QSEHVKhP9B43O+BLC/8QHKayP9Hs0ug2NcOvFTnB3EwlUxwXHlXUEi5uBzw
WKkFzeDuE1eSZCPaQfNfGzHWnqxUy8KBUF5uETszcCSvsikU0wZrYh6L8araUmxRAGNthtClbynw
nezeZCqzFIToEH5Ieylo8ju+NiQCx4kybHIWdDTqXmOQWLVGVM+nlTkLEUgDOnJK2UyF6SjQR8S9
k+ZAuTghn8/KKjoTMM/suQEhSsfGF8+VVw7kbUzcZ9O9LlAk9D0F29ZL+aRJnrNEUidvq+KXNrSI
V71tYmhzfeN/1tCGTHlY96fTFCXwTEIawWAMdUOTrrq8+eHrEii1lX1GiYfub+aeI+RC299Ck3sh
T5sa1+ZAFr2EsXogSTTuifNezvlIXXnaBP8Bp/bqPLwesum4yWqRMik8LqRoAe8vRroirEqUNS7n
wv+CCvt4WXiM1HciTPHaUbUPThhsjOLDBVWWEa0agV/MVZ1hRelMNXKPjwZ+KsC4H6B2vLurfsuA
88DxxJ0FtE8xBa4bYiNsNTpzHpAhsbupQPY8U+JoPSZZbzSfF0BxlZwen4jvoC6J8+LuGCu+Iuyy
0EaCVzIIbH2nxRuI+oBCvbYs5SiUHujLeP7XQr4z/4u3DKRDR8jBsOGLatdYaZP1PWFTfwEwRndN
t1tv770xarDGUD/9mFTnI64RnjMF+rakYOSAp+QwSLIv8eS3F+GGegTFG1VjREXEttkLtg0v7Ndd
Vfh2PwMlsPcVT8Yf88QJV378DwievIQjivs92Z25vl+j6KgyvjL4+bU+lUfdkMWSFwV85qUlJZg9
Xi+ehy1fsSJtxoKJbyTS+KUD+Leb6aQkJb2AontIidOjvrynY3iMmYyNyva2wU0kC3vEMtOfC3FD
IFOHFWhFqKKl/xFt9z4793cTCCHUFPwEzWTTA3yTohZhnAuFlVfD1LXUeEnVZdyNliS5KAXnwESu
L85VDFT3BU1e640W7LidLm8tFPpXWAe2IaoBCAetZD+u2JIq+r2hxTy8Pdnlljj3FJZij2sq0fWV
YpQTN05JfvlUc7i7jF7fnvoIs+PlxibRPm5AjznAUzOP02l0T19tK5loWO35FpZYEx6SLamXL5Fm
ss1eLXRMicZtE4vYAUWSZ2IvyJoeO7ExAubJGksm5fUin6wbTMTPC1zb8WY6KLqbCjtridRYWOkG
TXvVBVWQoG9NNdWVkvvdx3J2SHI/r0PHI+fizZvg3ugO39SHs+gXvEWD7kq38DkIlrIVpDHXJsdn
tnDdotAidthQqSa8Igzc9/ZyUShxsgEYxkB/xSLtDeElb1Nkdt6N/k6d8Nw9thWFWEIA5MGhEgxw
hkljmQyiT+su7zgcSbtD5U7nVmP3ejo1WIEp40UmjBoy3QEbozz13Q3zcNd5T6+Rk3wP4fusp375
gWSLM+PnnPfWT+AQDASW+IaZusIcoN30Uria3WbRB3VgiwpEZqebdL6Kx+ClhiNitpohLSYMiJdT
yqio42snDK6yjjInP5/nBQoO83+MarDf26w758hEAQP2x4G7Mnad3JW7himWJEXss7OHZPY10bBo
do2blM3mXWwCQWO2hwzbGKsaMm9R3qDHFgdDmtFWPAvGhSn4zyHGnlCzmJ5lsGt9TSmTVr4sBWWF
G3ORNwJ+5jfGEoPWhRXFVixBUv+fQa0Dh+GMgPaUR+CtMG57QS30j4WJgB/eh60X2RAlsZ99mdsb
DgTSdepc2DGHJUu4cqNsdduQ4bGJKkK4pgjsNdUV1JcO4M5/sjKvYF5wsRlb2vqb+4TZVDl8eKFl
fnqKfgjutfwEwp7Tgg2EAsLptfi2yRpfmokZjj6ZucTS9FP/jReLJ4aqW00y14Pa1Zgct6zvTPlL
1XlAplHjo+sDDfcw+napM2rbGDAt/E3TIFY3SM+BX/oOZnXdSUUJ1TsdTYqa+bkq/et20m4pCy5I
bYfB8BwifTvXKAJVOmNLaQ7XdAI4gnEJlJKSCqv6baiZGc3tc08RFACyTtj/hjQQrauyM7sxIsow
yWWIaMh6hREE8R0WLNAByfM1CplMimEdjIc3BE2Jems2t4M+D+L+LQ0Izmsg8T8mWT67csVT05hP
za26GYAvgbaM6UR+zdH9j5zBirM9LBhUHYkR/g5dmq6+qBjwiZgq/0OVsjgzpxFF3USbJBQx4gDD
QAKQi0reLBTVUv7MEPf/tFZL7601p8kMrDTZ8gR5YrKQePJfnyP7Amfo+jd68vT7wEJlfrKaEcuv
2b/7QD5L9p4FXmfdjUqmw67OKzd5/pHZU3NRg7+hBb77Z+cY94mNmeHEysAFRcqYDm3ijuNDX9Wy
3xoP9B19SBWtNJeGV5TpWu1UANQRdLpQe6F6/OhAps6NUzeEndTG2qpzHbT0qCcLDtNxrOZnSgEq
NMa47X5JPjOamxh/VgJxY1JQLbbpg31aLL9xTkBb+Ky9dPurPmskwjx7nNpJ1PKhzbtnkGUFFPEF
dmCJvpjRvvYt3aa2R9ejMgAMZUT/5Bmn/dmDeAjOPUDovdc90UPOT8V0KncJgo2f4AU5eSaoXyun
+hJV/K/3E6uVp3EQClPXPd6hPWOwbMRxN+0rGHBnvgQZO/nINP5CBvU7eGdofuh32JRqDd8NDuYT
LOO4hIDX2Q2aHKitkoYFTShnodN5mwOk5qhd+YGY1VAEJJldA+1BdJ8C3pmxxm8xEP7D7CAUY6n4
WqkSMEzy4cH3dUB9PlhvzW8cIptsb6/VyLDValdb/n/8HCTQgF2Uy4eeuRdmorerwKFtzAnYRpQ5
B4L6Swh3hlN5BAyAtg1RTkLE6wmsQTdAbHmWRG3EZweXCh2JJBJM9mv+t3vyvHMW/z+RSHl3Hh1Y
HeqLAzkIyzrgyILFFKs4X7vDR9dYNMioFxpMKbCaK0PwVoAZTbPu5vYiz+BXS6AH4oz0l87JbyNt
fla4GFP9MqOLnGdlV0bYWpePHbDNX2TaQ7/GW3thlJnTQPDdwJQIkGX2NekrrzJpXYKZZegMHrem
VJV82CGTtKhaIUmF55OxSNJqG8jU2PTug8q4U7bhWmAJRmfqIz5QQiTsJH3kilxb2XOn6WcG1AFP
bu83NjpbNpgFuitJsTSyngY1hGc7NQd4rjUqMroLAQm4+zP0rgzjPWCVamMczaww122QCYlITgUG
mfKV+3A9zCpJRHVvU2p3MfaDp7IOnRqp+2H6s9xA7cFPiKrPlWntrStKi5RaLllDlKZ9E+pV0WbP
81wadyvS1mhetYOjjvAQ7cdD+LQ1GYrwj+lhnx47ZLUif7rJ/kD+lEabeaNUUrqwsJkiINjcQoLf
Bjpp+xfjWzzDPeJeAFFtLX063BhvRb8yCUMqlU8BL5MePraTSDblDaKBS1EHpB4d4wMxjOBEhL+m
KowLpV0jIVD5FbkK8fAPjLfIKHAx/bBUCl0suFnbGvEH8IHCF3O5RY2tdSfY2CnhGknqdySg8KVY
6H6R+zY3T7Xq/IHJuFqYJDRilMmq9ssMmHA9RBpABn2Qh5884cvTdPpLwhtY7Ld8qxirQ+s1PfhC
aWJ8eFZX7YWOAfKulSXb3uj2EefoNMdH3P94FtV4lMxb4cO9HjGx7RIPiemEmI2rS3M2vHiGnmKe
V/drsboQ1yjtiAp2en4b2Gc+WbQMoDqOs5REwPlVo4x/HAiSKvS9ILPSIgZsm/LUrgmzkvqq5I5j
je8am7SZYBjQntH8f2u9QzaNjoqtte0AfBjNfY8XykMKzPDmVL3BGN2r7DNdBsTOfeSyVyElUM70
E5+RDZfqw+aELPxGbkiYTIXcohWMP6VgDDyYdtkh1Wr5OS/Q3DwDIHdMESaMbYeNOmWAmxHzV1gz
BzR8rvCVAjaTiO+4Qm0n07MvAIsXVQOhi4ILEqXoE6VSdyVPVd3pohjjcK/balI7SJ8YJk37Q2/i
j309kzV+0O7cpH75vtlj5en5pITaTt/tvSv57fuWTE+rqhYtAMoySW9jreCEOSbMf9RorNJpWygD
zjDhKjpEkW7i4jhFQKVVimH0xC0tECBALtRRFlkLYHt+jxLzqsdPK7+/xoQFL03exVSAHY/ggWbK
zuHA9wrmGdinRt5bgOFgKqdyV/kHZqdYg/n2Fwstv2NhtSSEiYVkql0N7vRcAXJZ8jMxnpgH/D4p
0J0Sj8Z1BpqqVGKBoKjGn0PkpIMva3Qs+t+pnwNCIiPl7eo/med/1MjjKdY6A9VEGSd6nGFgbk5p
B0GA8Fg1AP4qpqtbKRXbm9Z6tIyuLCn72nOGO5kq/e0HvJRwgkV+zCu1Ht8vHVIoLy3RC/6+CDuD
nrmYNjc3GY+1eIjNpgW/69IPM7FBsq/X+ulzWmvfgcWt1fIlr4hj/v6u3tYhnX4SEig1PmJhP10r
aeMoYmt3KRXljpCk+CZSvBv0x96nlopMyGX0iclkCvOY3mYnCro1Lj23lOWxX0b4zdDmJG8mcXbz
JTyD9zCBEKK+a01wFv5Mofr6M9yjRk+I2N5gF/xBDfV7Mm2eViz4AKVwmq8npaSJjYo3LKo1JJnE
jjmYoUbCtUe5nusmTaKAjs+Y3+LmXBnKIEMtFVMXhAPqoo8x1yqiR/3YS+C0fGmUx7pgW3M9GS6R
SVYjbKtT8SGCgyMCuZ1lKXrmAieyRMgFPUfw3L/ITu4L2APy+Mvd62rTXBu0XQ7/FzAnptOrpmpG
bJuDKQcWW59L3smp8x6jfSaeyop9wXsKsNpuR02d6+UpjDchyw4xdKT8FSI2sOzMoWjhzBTl90PG
VIC6LbSC6Nlhu7Vn6+49cLp3vKd+HjGPqzgPccwo10WbUqzqZ/HSLynntW1bNUxELiOyK4AAjKvA
Tm1xAWmM9jx1AFNxewT1j3NQcwgQH6aOE4Ah1ssmFe4vjwvvbu9scuOsNamsHGtTI8jEWF0eejmR
PT+HBP0g0qoeI35TQ/OT1GXMrGgMSn4T67CfWpnb7peQjJq3DPRZvw0Wgputb3dyv8o1064BsnhL
JO+t69TNo0pjZXCvWriSPqbftKHvdkQDxsolpFrznRc6jChqHwljQSBz6ALjbVHFLOP2YEhSTiLY
TLXRaRavD72p8H/hxS+vNE9I7EzG1mcoDzJ8R+3yRDNRGo3C6QhTeaIcgff/QFNWyHLwFAOYv8Il
tuHwvYlY3B40vtlfdJL5SP5lPKGYhisZ87BDZMpoRbM6kY84IKRC+fulTX3B8HpAi6V2I7Ev9kdO
84KF6qd4+lbSMv41+iZpalfGj87p6SYxGWEG8K9MOaT0YqpSR/z61NS+XqCtF/r7EW0fHGTov4F5
DM1d/6S4exD2S4OGCNKkL5Jg+4mkSYghRVACcRUmAPBG4Vck291PJw/l01qT1Hcwtqy5+FDTTzBb
oVxTiv7RC4mpAPCj2J8pIMPbf/rq0QhbCTao+03ybzZOEnDb8CBykp2DxzouPHPxfYlmD7JdN7gs
bY1oUgU1cw7ywMtveIbf8lm8Wsru8yxDOplrq9xcQ2nU8HnBCdIqYFbcfSHq0WM9ZnFFAITYFbX7
3J64R9TQurKqBt0+Vb3ml2QDgJR/WN+wSC/kyK/2RKvHbVXbcTubjESIge1ops3az7QBaI9FTqTl
dZHPSonsjeI3XNSATgN9rqqoUAdP90pxDRv4sYLT7Ulmhq2r2+98R87vL4MuEnBgB8aG8LnxpjqO
weeqWHcDra5FGF4XHSJQdRujgpmah0LXDHONdNYDM5DwYCFa9cvOwRglHHzK8EDnCU41c1PBSf7f
CMZgLDwzKSxbs+kd0aMK79HfSIav1jTUEZVL/t6vfAnimm413aNVrhhFxs6OGHoCii64yO4jv2so
tCt9ivgzguhX5i3Pc9IVwWJwOJgS19Jn4ufFY5/fVxnpoeR2g/D+oGNyh+2EFuL9mvOM+9TT+Jyn
edMGrefNLxE3mjXaNWGzQTsahDKCHnaTRP5WODVuni55IQlSbWMRlUx1i6zecGFL+6tfAWsfQncC
RUsP0UHIFvrWZeATAUhNwDxGyIbv/Zglh6NLmWq5Ep32zjICMGJBi/Bk45baT6kEkZoBEzEigzZ9
W1350KyiAasw6WzmyIVC59gjSLuaF//R35JriYZ9P1my59M7JocXSBf88n4adUcrG6xLT5EKXEDD
SGKcyD7jetQUYhyeVzEsKLuyILsi8kroGx0GSYmJJNCQZqlYwJ8cBumOjP1KKOKrxjsJ7eH3vzIA
UKQbvO0WNnf+8AEkE1xO/puytTPQGnyMSnnIX2C1DDgQCiCnAqI7y612VDPy9RJVKHr/14tStJ1F
cW5ljPAu0gYYxnPqVZEihs0TkUbXpLMt6lotQa3x4Y+oZ5g3duo6vLPGJMIBWgpHiSsjtMcMc7WT
ulQyt0kTBCvtbQncpQh5R4UZdUqGwgOBWpnIvh381ktSaO4+lVk828IM/c6+bKN7Hto+DHyin5RI
gYj2Beu+5eq4GMbkMzEvLupPNaPMoIoaVPpD8syOkMrKtQgBliiamUB39x4WIU9eojMMcEct+b8U
uFznCSkURKiFNB7OJqeeIS2rNrpkwIXaFI8p021byi0jRv/R8v0abd3yLOnY/fxokuuF5LOLyiN+
HfsQ/zqAJPogkfoVHEo5Po+NOXII8AMMcfnK7KNKr+FHXCF8NevW7oUqyuwITJOZUAIB2kS9EMWQ
jM0CSYTMuVRuvmOTuIDUWiglKQZdtAAhTWWoMZRc3s2IPGEx1NnxH4ZlD0eEZn5sxaH6Vi711ahh
ZJU9uiMzJAM6jirpwr437tAL/S4AeLsn4KXZEg9xHHLJ3PA0eKMtwPGphIJHWgJ0xVom39jwv7Bq
uxuUCixllBv8f9OmQlbc2xcUuxB1VHd6ACaytXv6vDDfF4mcstyCH5NHzleKUPttc2jzZZ+MiZ/x
usBCj+xxgRDTquiTJsHfZBH5yxJ4rsxtJ9efnFIOxGQPBlahxkgx+YStKwutRg+cN5zlHe0+jJRW
SDHbg2BTq5Uigth+iPErlapxX5IH3oBD0SdNvedpXfnCMXoEvPCTDi1c2hifUPHPYoNktPFe+cEd
AieYCTKCBqQqrgyl56Ep2wyF7oKCBoAIp+1vq3E8j6aSHVvRkdJSVI5n9KFeGelE/HzzMHXXRbG5
fZHwFRuJTun1XHlZfgyPm2XDoCEipNh+gnFbZTXujPrX+sgBC9OLJatlTaNhErxn24MR0Z4iRw/L
jpLxweMi1pl1iv65QJsvUG6CQfWha1o1RSOMP66y5zQv9OFcTgZtKL9i26TEeAmw7Qzd1BfPnByL
C8F/V7dWPz0Jbp4ncCRzBm817qWPNpRt8sTRNy0mPXoI8pI+rE9VFbWxI0xAOQHtMH5pTEce11PS
zctnAeBG62KLU4dwW+BTHrrrgWQA7uPp+UnT+ejEJAlLeI2KXblnrjGJbNc1tlNMNax/Eymvybhq
rtE6/JoNx5PwbEra8W8WlKoEExTTZqDK+rw/DNrN6fymeTMc/MhuA3DiIZwPMHdcnu91Cdblmvhd
A+XuOL0pSkRuRqf0sqqxNxs4mJRMe3uEuADcXiYVU7lYg8hvMji8Z3gVbpnppjQM9HSDn+8IASt0
btWxlckTNCEGGkZLDBvcRDpdAmWer5PHc8Secn4BfXmTvd+txylqrztjDfySWwF0PVKzK7gdlTy4
u5JOW0gpeHVCmF+c/rxehBOGzPtUgi7WnmIMUhNQoFPSWNdiCLma/QCWb/T+n+74EZ0G2jLWmYJ9
2IyTqFs96N+mniS1dJLDfhhmQKfXy/qD+X6g4yiu3mB2OQ6akbG5ArUlPBYM3opBClI1Qh5jAty9
ESYpx3k7g5GkKkUHJyv0OVkppJVjQit/c6g/6rORu6wc66z80A3y9SQSSTLe+MVm29Kfd3yVX4ZN
o9uz5sfAq9nDvYMwcueSU++ddIQmvrrNWR+PQBuRXvWtKpCKHTyvsYHgA1kiyPdek4eq5bbjfX2/
yMJ1l+EDCOL+Luwgq/bHLv4S2vX8ekG7C3OgiNYZwEVlneH0xC8Q/vy5T//3mUnww6kiEBPVUsAO
obphDNe39DXYNC866P1dIv/Gr4SihqUv8UeyAkOs6g4XAOc3ZgEBtr5UiF44vaw1L+W79v9p81uQ
9gFbjp51EwviBWoHxN5w0T6bHfwHZt2DWHBRKJ+HxNwELp2g9UHbrfsvE1R9SQCYCZ1Lz5W5d7NV
6TpayjLhzLR854ZcmmJ1xrXv/FiSytl4BVUJNYRAAw9gsOcQHHICJVAE2uDuQdcu9vlVCGVXaT1f
4FhZpIUTlyvwbCrE9RjlFZNNEvx6fwWLlrIMZ7zhHQuhAJLZLgcVBZT6mdfLjrjs8t8Is1j9ak8Q
aX6FqGI8ns86v96cMrVobgkpU9WAd9fRKMorXVx+secP0M74EVMXHeqZs5U32uVhQia2mZsj+X2h
CgqFA6MmG+OXFL/g+GSihItQELWoeoGN6DYwhQMHIb6w50MJ39qoHqaw+CfjTmNyx6lNWQin/YQc
vXAgvZjG0+aWfIIz+ZZDC79eeoMER59I6izPVZV5n55Qs9Kcbf53gUKbEhtLdnksusuL18ox4KfG
ts0AHFlWI5aCjTMUKtzbAzsw4RXMu7+/LYArY8Fz4/SVThlTGedoVRp3L++GvZNVA6EKUr1trccO
mDAzmyZhP1F1vkcsM1RzBwPbcYeL5TBOqYkx5OBKjNRkT9uOnknlmEvQH6S+DoISDBnG6s6bKGfN
A1rlsAd5XbdH20fsLbHdqlN9E14Fhb92/CgZNBDpe1nVdyaicXnXS9j2N3LjTeMORcEiXlt/aCh1
+dKC0VQ6E2DFgflRw1nlNp/pF5YaRB18x/tlY8W+a1jmBgqjxBFiDEHpk3uj7XesVYxUHlIw62wC
ELoRMiL8DyK6yTKpMp4tKtlu2hwS+1ZFlbnhPgpuFghiWLd2C3pxCuQ7PK/D+W3vtBY+XOf+QNih
rbIKfngKkcrCfOECGf+lLjWrG2F7HsEXmC35Rxv6VrPWAJG2BY9OQO8oZnmYpRmDYek66uyknKt6
GR0UtyydD+Vgh+AWQ5Hs4xoNen3dD99U11SF32Jvsg/mP+BjP3AyUzVMsnLfK/hihKRvggRHFqhK
OOuvRVIHMmylfITZ9xqHHeWJ1FhzbtLUYMRz0LX2UHqxQbTybHzqXkVQwhvnAKnl5BQ5llS/pTLW
Z8UiDfJ6vke1lYE8Gt0SowiizFXZK70C44YUZnTnzehGwJkRqkxOsdzKDSMUH0nFFQvAkZ+dFuBH
cqUklUKcqCiJPLndxGccpjLQVro8/ynKf9KtutwE8+da4KtXRTrjU1dfYzp2w3R8Zs0awrWhDTSs
vgb72Utp5la1lrbpk2gb47LQWODIgmSfdme6uYo2u+Xf8wUth2ncIeWMeJVbajitRUVH1EQgaC/r
znH5Ju0F6ORAeYul70UlB6KIq7BkslPriQPwnxDno0mTeDXnVuawApMH9Tu64S6sdnH2f4IZpLDV
jcPnmZVG8iTbIr3QhVpXJ7ZpYbLg5L7R8RI5l+26lNuCTGo7eaooIuYsqO0Mqmd58wqHchWnfDOV
1HaZOZsOaUte1dsmy9JOWBpNpjM10PpdOo2Q88fpXcJ75yBBjh8WLPLMhkD03fVRQa4xm2dfhvWj
NxILP0FQbs7WZoWCnZvhka5lZzz1KBHGJNWuaenF85gECqtqrhPeOQIKEJknv2SJOnn0KrUNbgh8
aweC/jCEzVLTL9nkqEGYBCKXk8pt1Ej0BJtuEYb4nP3r0Dyz6b4ZRyUUXcdQ+YCrYZzvVIc7dI0Q
ye8Te1RN0ZXTWQbD7H+70bJmJani2Nunh+N2v0zJL4PJBvjKsN8/FjI0b2iZuXGzS2ZcyKhm77Q9
M+n8qVVHOqwhivOvJzmh4v2yrOQWCmV/wIEX5MV77jIJ5PDnSHIRZFBuYQk1bvhmGi/Nky+hYN+o
PHTg7ta9YS+YYTqz/1w+ytdnG2wLM7hxQZBqaM3zUMorbGqbgPP9cS3YYyn1ryp5cyGcH1SVjD1x
xLcH5sDNgi+q0Pfgj6VuUxe4trLi2Nz68HRMQAPC+HjtWWpoiL3jN3eOU9VBlG/FXlBgfHBIM7Od
7JXJ24UbggtJ2VoavPWVasqHzApCM2PmkMRrdbeackz4HDHHWXfGWjEbpQUKE/pJQCC6XuDMqdZs
yiVTaK21oN8KaaxrSmlDa2N3W3NHXxXyqsCKpU43CzS8EBEj0UtRTHs6eB+47YB+LHPaNSQYRvIL
esF3KhsLWlU9VSTMJlKeVeGTH2pZfU62Bcw8f1A4sHV8Ac0TQ9k4CGv4uPvHrqAM6IHezLwGKiyn
3sTNW4PjaQcwiuBVLnzvr33lEYqBv39Pll8b9DL8DlXO/a0zUs+O30o2jme4/ML+oRloDc7feAmP
czIN4EX/bbg4GG8coziQLmT7OjyjpDehDQ3wwVct1xz+jzNg7I1oqEUmW3j/lwhjYjDd75MQGh21
1CVaGnMaxckAuf4jqLqYE8Scjg7EAleNR0D4BGjfHX34lgd0ZbFXMT+KUHwqkwe4lR7r5nqnVSWX
1v9WrkApO1NW2Z1EdNaNNlDy7UhjOvh5EAAVOl6SQ0YpdRVNYI9TNmoPNJ2mTig6qIvfcfadp/Rk
Scw25av3nnpuzs21CxZilDqhBeTPICIaCCJHZzPBnS67sDUAtZNpYJ72qZnw0NHcbgBjjOK/R3iN
/eYWnqAfuvwzWdYrKdO5vGo21g3Qaulw+LJy50y/K0SWiRc+i0GMD220gQJlHtPUO0mzWFd3O4SK
6icXycRsXHatLGsS0q1EiwB8j4ZUZmRmXBX5MH/29/M4B3k7yubvr5Eoe0b5116THRooDaCJTJFY
8wZ7P16IjygHxyVYlAuivKq9Nm25J/dOGkVDHVlUd8gTNXWn8KJpgA9is1zKoiY8UyQ2VVl0EkIL
oVY0XnvbB/ucdWiOc+J1kpKIRrmfdlcxgYtbIOHIyv/s1RIwhV8w2hG/mcbGNIJxTMktZBuiP38n
YWHJL/OPco/fOpVVM/1z66sgmj/5L0JLPNf01s5sZBU1olGIQFpFR+yjD4yUe5sPlonP4nerNuAh
DxY5pGmRnYQfzMxlTVd6aAlShYd2zsyjjA1KLxLwd9FjsbsjWJGYsWNHE+A9OmMKGZaJFgBqcoFY
HtrGOvBhdBTrMBl83rnQSwTIJ9QCrMLhrriR1NPN+trk84LvnN/Y/9PtNBEVifSqc+W3Vi2vqlki
ik+baEKS+dv6k/7DTU6If2ueq4jX1pn4KxGSyXOpdgpqQVv6jdUC8gahnk0sZaN1yrqDwvCisXkj
afdM4zRlEFqwaEjZnKh2jjObr6H82jvG8bmjSQ6PP0RZ5D4SINPph7RQ3FfpxzoKLrDyXDeULRZV
EXTA6N+G1ezTBJvzQ1xnQJ/stw8W/voXLLiOENBbBR3n0RS21x5nIa1U/a+S4zsjpAKNpcL5ikB5
v3hCFwY6ROj8/ln86s4jCaQ8nme9RNgAyh7P2aYEju7uOpuFPMooPr2pieRUcSsBBWWZVdHUrG6G
vq2a5zYFXVw/fQIMV280eQ1OdvSiK0uAvxkFCpQy9AEeajrxlOq8p0ehVXzUU6UDBrHOW3IaJP/H
1RC9XUTHbTu3vRXvyXNzFMPMBL40jm6Cr9AwkvEyuF/7/9l3NpnX8to/67yvi0cVjqk/Sj79eKug
LuXneMdwfnlZzCwVQYzbO0qC7ckzJe9RcIJqzsbQc640VHkXWwDn1IQM81xh0tZlWiNon3LtOS/t
/2i3REE4sTTJvWpsYP9fpqzP1aCpIUdk/L72k9VvcA98mgoLRVJuDXNaZn+mJxTBNql8yU7c7eIu
raL65+FL1mBWLOU+JXvkyFwcgTNAiC8IgKbu2XpW7UvL7JYuxeY7PjUL3ZCgEjMNxVlrSyjjEnVX
LNANusjiYvcQFME1IwHIT0LT5eR15/+7CS34Jt189zuI14lHLmSa5iIT7DKWs9bDN5kdeU2FZDMR
wmZHT7gaqpmLrefDRaaXfckapdaHko5AFiVRWuq7LsdSFN4SO+8h+MjonFlu/kymVpZBZPTah0W2
YGIsa/KEWmVs+YSL2bpXEtEJsGH56Q5myJbYAiHocvtAagryWlr2PQXZoQDkYYXPvpoZU2tTy87Z
mA3lKmtajn56OVBp8nhinLniKMzzVKhdIPsCtJWDl96vuU3GlskkUzZLm44OpcWU/ZAB+Tyl4Awp
w6Vom5kmJTFaSZjpZA7Dztl9GY0mz+7NXEu28fzFPWL2GFfh2b8ZB7TEhXj5zSOf7zeB05uAiazk
BymakpbPxv+KFhRuISVTBtCPQFPBMAT2f9UKXc0QPhdAknt8A1lH4pR7/AQexAWPIDpnVhrkDrc0
oVwxdAYAEwy9gmYxFNxvGX6YW4JOQpDhgecvvAjbn9Z3i0XKq+jvKFJ89SrF/4hOyIw27ynJ5xqd
OXypCYffR5QdcrQwKOM8rUDTHWJUi8DR+oGRLfx8XnMSXpz08VrRMi10Yru+w9BLlFrJWreBNF5V
auADpxm0lrSevkU9LB1p1wMBCwVGpBt0u8TTcTqAZcxsCYyxsEk1F0GphMv+qllr3jxRTfFM2stL
bdO2CKdeRjZ6BM6uc/7v7/xqvT91iHfPFadgfQ5cDsvRO4y0L5jMCq2kphBNwYp/qA9V+LjGrVXo
ENuI3L6LIB1fvzXmgmJ6X6RD1LFF/qCSwCF2SioMxvomif/R814u1Lbq9cbiilK6bYxGqLueLD6L
FbesuMjyC7c+vmU4SBSmf3t5WbYEovwzyywrw2tFr6cq7xENGtUeuRU6dPiAJWeCgOfDtRYc7OhG
16ExAloVbQwulrfLoml/7gtlWXQtTVcHoCuVM5ojnHzjuytGH/zyXCvmLmP7NXuNSvIxaYLdMXeJ
892yxjo5wroYC0iLqrytGoN5Zti9/2Ifa2CzVh4wB/EtLJF23HJfEXNIssA6AuwAAoPP5WPNuADY
gWaJdeQGXVzLwm1+OUVQmLSQ0U/CWUSEweqCYTANnME1NEoIdklbHPy2r+BMXFzMB7PFgEMLfUbL
Jn1N8uEEKnS6VXkxJyjyyn9KXgcM2KORfBXjt438gkR3mqLRR+zJmGw3QmLA3NwktN8YTGHF2/qz
RUyVI7PE487Juy4jGsCNTtB27SKJddi96W9WZjAmPkqUwx2Lh7mhibHOnauYZNdA/onlK9E/jmvn
/F7/+T6m6R8D0bymdqU5JeEYs9ZiRH0UmLM2yg4vFios0V8dGaZRbRKrDOplInUQ2ycVYzuhvotT
3JBJih081TR3ZXw3X3v5sv6TdWRYU5inXOLTRLtoxP5q6kP82Hy4PEprN7hhhZYSq43JekxuoeMX
c5C9ak84Hz0wRxVcFdwf5ZnzCFI0vNFESiahDfeKHYAHDh5DclNnSNyzVDuPMeqikGeQOzHM9BEG
MqgXB8YMySfi/wVioot0jfWTLKqpqUrYXjj0TZID3VZExVJKSuKjjTf6M++tGkSNBk1uUIT5tYPN
KgfOg3rTScRBDFC0YZLVJ31YC1VlTzscNLLdeFTVEZtC8OK7z8lWro88O8gb9MByBQTOJ6ZlcL07
nx2U7bKqHNqCAZSx7wIRZ43ZJId1gMYLN14ghTc2ieY8nvpXLhhs0gXv0PNNKkBlsfxx8/p/mJfJ
DGXhEEXPJ/a/Q2exMQ2GJj00HJnby21ANpwg4tTvCG21a7lBgWn2E0H3g/MRRKgesA7numQz6BBW
kgKt5onb1SgW5f/1iQBs9vDpRvPMQcrnPXmsN1whhBwjjl7FHnmBJjyaktL8XpvUTM3BTSyHTn/p
11Fdbjxyay4ZmzK3irzJYrd/NN+mLaDf41Y/X1ufrb+R7ZfWgbAi54c6Mao56SSmnB4ahpiZhwIQ
rOWoyPgKmPlOILBFM0sv+3SGrB3iIbn6LJUKdddFVqG6vjZwa8Y7+NnAmxEL736Dmwr3mbFG4LCo
gaKE1va26tshMxOWkxzBFRc5X3JG2TNLsPgj5jmO9Hp6MEfGIcDhSw3u5tO7iiWKSUDDELOoMPdu
YZ5pUCWeKfTgnUFIbQ57NWPVfimpg4Mjn7iSg5TdgmkVPVPsUyG5hLgS6kN+3DtJhVbISdjT4DZG
9yDYYPX0h+UjkDKYqNeb+ypXnIW+nZQcoMWl6+wd7QzltXlFoGiJAQyjF+McQ6pYxGQBedlLYcBd
VEvq5FrSDkpxFBWVaI1hDbzhbNC1ZygEBYeEEvZNknCBupXopKMfCUWsRg+Bxh3qgcFyUaUannj3
JubESDd8d4zPtF1fX+Qm0eHlB+qxkD+0rlLZyuRBxuQxaDkSWEMRK+RIk79Anu0W9EHAmLaYtBs7
48w8ZwTzXYdqeOt2qhAiiZxtUKb2AwAGpllzsYq2YXNBTz5UGqy0HKNt48bFVs1iPF8ZGXXjbHS2
1x5t7Q4aGFuSRzyFizELH80DQUGXFGmXzpZblKV8Bhje9gAZ2CUUuDzEvsT5+ki/2FuhCq/YYZEs
scRyKMyziCNMPykelKlMs5V0oJrd1sxXByCYz+2NHn1sKP8XuwJ4Jdul1y7iOrMUb+o/jvkfVq6O
cxYmlKxdYExpNwMKySYISseOW1gAu/J97iJkhaQG9SNXn77nhN+9tSY/2gjbxKZFuBEuJV2G86iH
rQImhNHEBGSj3FxgQSIlbz1feTHrI9E7SgB97WeTn9JV/HUgvHkTYIkDyJTkgE7WWMFswAiXGwjX
8aMfuLO4NGeOTuC3cfIwsThFP2JMI8DFlAwSkOLJ2XSYsblz0kWXXfVbeGoeSPkvY8Hy7I473bCx
DBvg+femyTEoZ1EC140XumTYGorrpoFz8gH9UTkJxl4fN/yMAhjrJi/TjAWRq9jd54OC1KGowMKo
SdhuZoeCSF2AkNo1FGDtRik+VkeFc7DMOt51tNiY6W18eyUO8Ae35cCPYfH+i5lZW6VrCc79lUSA
B6+lpVttyIlhfE+4BkCtfI3nHWQUp5hNTNnu9q/Bl4neaPKOCxXm7XWp5JI/S4QTTWy/SuE6DwTt
3m3QtL0xRGACtcoUyEWKvSd7YFafpiMv8/F94QRoqTW/dvneLIMobimonDOmY8edxSWE+4061ATZ
xxlyPwC3k9GDatwVO/lv8nmrJE6Rc1k4vwcYpESQP4/4da8tfwcIB+QR9L4xVCuJr+FgXP1W3F9S
tJ29UGftRueCUG0370cyoHlCgsa5elhD9CLDR5nkdaAdtXJFIRJ9ku1x1Shy8OWfzRQN0D3syT7M
lNNglmCX+1v63HGWtn7E+A1mOFxQsPfzz4xNfaRAJyA8EIf2J3O1zNNalcHbjtBgGSBSZ0Y/Ynez
ZXufGIuu8neQKCnXcYETbByzNlopTHdJoYy9fQoY81k3OX74BAaUqJD6+IZjrpfN8yXsMdV9sghG
o+lIqrseGT2iNs1cgMWMYn5dQjF6e7qs0GpLL1qLiW6vuH6IOwssKF8eH2qJoqQpFIAoiNbp5Dgc
P+ElMGU4rZvTyI2PHYr0PdaNETwl1wYOyO/46nDvoyldiWpwVFG1Zu6+uN594poHcgctlTNxd/f8
1qNF5BvVnEKtNqiDK7n3cpRk9Mv4DDBXA/bezbEyAfi0S7hzYgpbGbL6YquPukEqb1AxeyiFZhvi
YUIYUEYSKT1KNLQLxL6Mzk7gT7WxoQ2B/jLLAXObS90/c03IAYW/Ob8hk2lo9o8K7nrknxxfe5ZF
GiQDCoWOPlNpOo5CIre+mQp/b+039P5EA4RtXcaLBhcDV0tfrkCyrewiOQbDPW2tAvd/c7HO0KjE
CcCLCBrNlVYlxJvsZtBPVTk+iTJAdo9SLVJ6w6CQR3UohEbIKvQEKq4Uh8nKmne3J/vNYR8FkFYR
KaTZV4dxaz5bCdfGJ6s7Z9IAWQK/P5eR5lZ/9f/+wE+3lPAFVlu/qlkTETVWf7PEjEslstG31IzL
K/L2RZyAjVaErc04UXPk9OLyVy00KKEJT11ltf4Iq/l44CpJ1DOKCfnyHJopdw7iCQZ2mOUTnE48
ZGigyP6Ib0xOo4DqQ8wTbqcWqz17y3h+bdjJVqKrSXx7+R/82rohEtoUFNvuJCw6v+nrmxOObRCF
pukNwwvMSy1ASP5ju5c4H8qDvNRn5mX9wjYKJVDuabn0++y8Xdt3MkF1HTgDI2bTLn81GJXSB5hM
wtgk9OGas3sTtIm0CTdWOTjDhTUEmOG1OMVLgCqj8z0qzkKULN52BTj81AbTJfGRjdxo+Esw9ilr
999hkStT9ecVdgISm85eMySG/GT6GSoTQGxECKdzFfpU/WMo3QjXq9sppSIQA+4Pm4Idx28NYWY2
rIYkL9F0IbLDlTwBdQBoVOeSGkVLxrgGxNfdkJsFc2F+WDaDLzRJ9zC03e78Ff8vzUV39P/gywCg
O9C8gp9wzBSR4/If24S4qYrGd82rlbS4QiATgTffgnc8gmcB4bTBRCaxWvlTXflnXEevdR0d8R1v
k2as6LAwnPSWYH5NU1qOYsWFCoXzUVqGRWQGbLyVeetmbKfFafDzuICo9TlIQzCibxF8DATazGKn
ltu853H/ZTmDI/zCOK3WJm8/r3rlCdlTmRqdecFHtLRmkk6ih8yjnOedhEfVz8SJf/pvQ1s31WZ0
1wGClkskxSFGDWPpbPy7x3i7E4qH3hgxFJa4hbPtuTW7zmhDX6ECPKhmuMAfvXk2lzi7T0g3be9f
WFKdii+vtqklp8eE5H+h7u6+YnyrQPv8f3hn+C9qsnx6HnwAmjj0O7sMehMmaaDJ5gy84MN/bryv
/rR1ydD3pVC0XdEsVj76IJmuuUp87Ie/iJ1ZSLjz2/K1tv15f81vYl2qHE30N8n/NiQVYNNX9h1N
YE1wvT8fc+CrOkk9KOpxB3FRZ0W4maPN3V8fZkbgH/CutpSuipoR2/1v4r0SyNmyVgZIEi2B5hy+
khHiD1lh/Ea0HI5RE/+TM7e7sOvqBOHCgdLgg+gEjUiHJ35pGgJ8xgoo3VY+wG6IDjYN+SuXevoF
ul2c9xiJABQ9a3+aqG55KC0bRaTn6hfTXnvxr9DADf8BHrIXw+eX33PXYALYnbmdbDGiWM/nSL2I
pl4t8mx13MxrQUSp3rMAdDFrvI0nQ63Ii535v9qsdbDWcA6+j1IF4CFYIzen18JPIBAOvlEQp4b9
GOsMOKzwtHUZjiy53XtROqY+2IfVW65/FX9MgBEZToLEkbFr3yKpBg2rLLIB1P+F8P0akujOi5eL
uA6Hxzdy5zC1lcP8LFQ56FWtE01uHmQEY3AlWdPWMY2uBWWGSGfO8KOtmY1uRE/LYBou4SaSAfR6
nMe0NHgNImwH528ekOyr/8bJuKIcz9WzNQszawH1o4e2tXn5CM+wiFHMXn5OeDOTQDbBJ+r+VbXN
nsXSw7Y2Qxeb0CGVGtNCBols8Co/Jnet11FoQh35jl0tz1zFUOkj4rXGws5SjZ90eMZlgvpKFkP0
tw26rTjqr3+8tkvZkU3AMCRFQnPDK5l6WL7CT7D61SRBmhA9DA+KT2WrL3hkIj65FfbekAVqOzaE
DcaInrIf35K7THbWxT89Dweq25ooqjNij+HOT+Dz3x8z+WPirooOwUnrwOUPbGzEqZa0JTlzn9EJ
9sj5hVK0CUqgjRFxtpABzyYeuvlkCn6XFcbWMM82W8u6u2VP6a6jHjdVZaa3lG7u6bmoXZJUZzUv
ZDHtm6zOK/WLHiloIkulDF9XPWXIDSSNGuflx9yRs1NXvEa+0Tw8H3lqqvAj9RcZoeRrLvsjukKJ
9BaaVIda+y4d0+mzipAdCYm0oAeqbAIPY9iNEVBKAfCtpSrfkDh4bJjj7dnzzypJ27SIqGySVQB7
J1e6Jj+8f4SuUWyZkK0y5EyZMfTrJZCEs3kLxMuoTpGeO0d2e/wFr3RdUA4HBNT3PEfdtZN745h2
hzLvAJvTr5EPwVO+MhBvW3eccUljyqmspXSaWKszNEMwiFd8LYlHMILnfcNwoDLNKd/OG7GmYATY
ZOe6r4IKtgdxKoK1PYD/VlXMBsQvLoWBT0Rel+0YZJ+DyMlS46cbPQc74KseRQ2F/Jga0s9eSFms
QsbwEi+WKG0dLNmjmn3gJ8lfKLXKW2BLl5M5OAcmxIuCfBWNZv1bBKVX98xNl2SHtjkEIq6vviYj
gQIw0GLf2JRrfVChH2gz+HDJMvUccTSSLGpr1SbRP8aFXpuHJaejodo5ibcfGyrHL6pcNfIfz/k2
PfJr93If+gpQ0dR2nKtshHXAn5IjttDJWohK3tSEu2qXS44l7DRfhAAFjd3GFtemF9uinyA0z17l
oZZPdkGFzF+PO2Xd8zCx7G0/TVQGPX0YuHrTWxUs0UTdjAbdi7M4/Y36ZZf1Cm5dWCrIpV3Q/i0T
dsEgNn3iueknNZ1reQA/OavTyftHzctfSHb9Rts59yqG2RJMImZYaHESagusm5p9F8Plfth+3rmI
jOc1PgH6gQzO01d65Gl6JeKauUNobHDD7Q0tIgN7nb0qlKqL1uaIlwawuNkFEgDqwJTRLc/LV8JX
f3fKNRGZomHsNjqQUne+YyahAL3UyZ+3Vq8/RAzLLG+88awCV8LK/FnE0fA/inLm9EMvtNFBLdvx
LzPohfSFocUFMYRWXMg/BfQ0wWQDg240J5rpQGGYtba8GHv+Q49qaZGHe+5Bz6ZJDvMc+ufDQu9R
p4vDNnNMc/WHxzBohblELurT/C198v9pYfiPVYiOYl/MtoLGcpOPTPp2dygMyva4b8LVz+L1O6PF
KPcHKn1DfyBcw7+ZsQXGs+gmc1ZlnHtdAJEXEwtFBYI5bJX4kBGaDUYuX1zRrIKyCvQyXfIt5jyL
HG5fecXFsSOw7PS7heBkz63p/zg0/X1fnVUtDQS3pFfcSybPaCt5/8UXp3sYJXJ77McVx05Zj6AV
3sp2l2jOXclaFakuPcvbhjRb/zqowASiesiSCw/Yt365zywq9yXprTknHMWPCRfmEJ93seXB3BIb
vLaz1l0upVo4m8/nKiI0vgLFe+4nGnDvaHFk/zZgkwMkUokeiDgTCBI+qtdZLYVdFZ0cvZ0ysexs
XMsD5/11uqfDOS9nDrS5yJFhGhvKBegOYBpKeQKp7emFAEgSxPrMt1dSc1HdiYUBCJWaI6asojS+
/2+Kxv6eIKfapD4QCif1h4QWcN6JtU2vmmq6ZVrX35fg5bz7l0oiBnGG+4bkGUE6Xzkc+Gn5ucB9
G/teaYAkPGTLafxItwsLNSgwTQ6cz8HnqJZAYqqWQ5L2aQy39QCK1PF7poFFcxQ4LmWxaEUmRsog
txXNimcMOAtisAHrwxS385qu3vL5oQkIbkQrnTgfIW9573xOZxwmKkBJdlmj+CD3d7hh00TNEdtj
w7yMqDuYXdrNQ7NkcO38T456mVaq81Yq5LKmkBebAsgMOkuEzdzTr8TuNkJfhAvfKj7gjLlubqLv
D7hL5HVV8JJEyqyRE0Cxei99G6HjiMbYsaVu3fIVu+Go/RvELRQjD5WdwSlgQOYrbYtjYi/Tx/Cc
Yu/OXclHwWfTa5KXNnsZIDYWtKAolM8HlXTbDkgJx/qnMDT4xROlLFvRQ4x3VfX2iUEbkEydFXz2
HMr4Y8/AgXcgJuCsXTFE21lyEr9rJ1UFFczr5DLUoZYcp6PKHEOZco4GWMTGrQd8OB29gBTlWrPT
CKXhsOPQ8bCZVKX3B150a2JmUzFRXJLiFi9B0vZUs/h8/U+yXtUODVzwlGyReFX7Uigopg4JUtiz
be+TQ65JVVrtiFj2ugq4Kv2Bql/k2kGPTMAESQ1hJglBZesnGvXacXeQhJGdru+KW4ZofU5X4gV8
eIMLW2Lea1mc/fZfbeBmnfejBd9xjg8hAaRKzI5Ik4hLE6nnUxxwlT7qwi2s2oavwR0pryXkQJIc
jtAE8WRamAB9oywLa8yGUZtekd+XPwFmcZvF1ttucdIb4r5NQtcZ3yeZ3Kd/Nuiywvns5Q8yoa9w
tJSZcpRPfh59Um//QP4Ng+VXvtNieDaXTjlFt0UDd/X8oEE5tXd3pOU7xCAAOQYZuBn/U5saqm4w
6/ULXXLhafTqBRmYOiSGI2NmThoJ+Rn+Y0OJuJc7iwMIb2OzrHXhAkk3b/rYq9kKhywm5ni/x9FY
csKnJFRdtZV0GX4Lhjim4hBXHUT256mHiCu+H+NF5l/yzt+/2dycHjMTKwYiJe/dzt76soL9YD4F
HHvcELrvFpy+nFTAwxFLW8v1cFGp2IEMzjBj1LyJ1pLJOqN+KvL+knwQCsJ7A8KB0HcCQ7vos78G
PXnnAVLlrywhnfGa57CX9r75jrQLnbN0zbJwOCvHY9CYSWI1aIx3BUZ7xRmbj/xIQFZTNNmuPWoC
tjRnGAwBl+1LR/2408Wkl+YBLkHnVKrkA7dzHyLtV4JrdghMPYD7q8ELUdH61b5eS+CEUiG4EEC3
Fvw3Zr/NL0USH8ip0NADI486lBYlEEQwMz0zo2KUxbQPMYwE1tMMRID87alYonLBYy39oNmGs/Xi
EE8PVUgCe8Cbf3XZ6hpVTMKZpOnq7K0rxWb4NL17Z+VhM8w31AvIgLfd5ac78uZ/H6iuxYGegvsp
i4RbNLNWY5wTjG7snDcA0rznHts2ttoQv/JstGYTSmFVYQr3kp/WcWxsgMbf3iYXXXkkeDA+lBUA
H+GQSHVdl6Lp0F4gzUE5yr1b3JjFe9jnloWYXkKl2AWIueMNaqDVbAIjiZLsIFmZLvtt0BNQh8l4
IQFUXRmUq8mwwMGAdTn7kwhgyjoJGyg2aAwpjfnt2HzU4lsEvFNpG03v/FmPGCjOmWn3dn8pymSo
u3hTwznSkrwxhb511DqIG8aYLgZNVF9BFHjZmVfU6brseMAV4htJCxHoDvRCo/ZHvdhNHmEMiuJC
+i5GEkcKp9YHLIxNTJeLCasDyoxb2tm/qKCwuBWdSVXk/xTOjd2N+Hsj8a98s9fYKx+/+fRU/XeB
Rl1/BXwr/7V8xaGXit0cOjIVBg2ZkG0r8KJdRqN946eZh5WGf4JdQZe3XFzOkd7j1l3Q87/CLlSG
5ajXwHVbjz8tIsPsWKZzL/El9+Vrfe4XpiQtKS8QTXIYexlLKwekDhcPTX4rSEKy9wZ5bzK9Dejy
KTK9qAIphZ0rhIk6QKSj11+bczQmDUbppukVSqkPexpKLRUH93I++KP+lABmmjfhGV/deptu0JQT
zM6XC2eioBzxSNadn24HXmwQ9yiDPnVjsKew75XKALqsHKDUqgLkcjkJaNjSAfjdCAzdndq+I7tw
Il1Q2meAeDz4D7rXPjr+JGVlNFncozRyS1NetXQKUt6NrsrvyotwbxO+8NA58wVgr/DCjJyTb0ms
WahlfzNydvwu5nnsaq3dztcARzrEsvc5hk4hqQ2Co3ViOI4D3lWpKP8aDvAAbWsxr6O6GiNCh03W
k70pvYNIb9ZSN0yjs2TOfQsZT4W/qskpIb5A/NsqUu80RU1Q/FEQlmcL05I2zeocPPZTaOQFjE+4
3kAPHSkvxJPX5L0ZhY3UCU8b5qx+GHONFyLMl3YFQI8/mGFfPkKHKUe0mHvmnIBiY0GKZ8RqXWTZ
3Yxd3j5e+XW18vXSKZbATPawXdKF3pHEOZozNNXBiF6jfj7NifBYPDsdZBRY3uPik77YR2tAZmVb
tyPyyKq6zlkGn4cR1WZB8/by2/5SzJIXp07um4yQvxp1ws4JJyaPS3zdsgFqsKVUorWroqH7RGHj
gXesCPb9kB8K3PY57hyybBDFsFQoeb2wosAYN6TzjqzEf/Q8BAU4Rob7E7P6iazFupgzT3y+Pg2j
NyQy7zu2yl90n6SSn1O0ZmJlFq6R7yEvVxDZdC0Iw7cO1qTDgKnMX+ZkF2ROFwP/yFSalrPkdJMT
g+fvcu+3pA6t+6A85zlLtzhIbE7MpnHzopJXx+20zuZs6AkQL9H+BHrKfJafv1I67zQo+LI9T+10
KszSKVS2fpKB8ALzMJuZWNvQqoYU9CCz84ye6NZpoolxfNC1Ufy4lMqVM/lj8lGiftAss/3k/NPk
sH95yaktRv6Xn3+jkhDlwDrTIRth6oHdYYe4V4jxO9GqpobdJl09+i2Pw/YoDKrgCnbVJC40zvby
c9DlX9KTgZYv7Oeop3KLtsCurYTZA4GYjYTmKHKLLlWd+EVU9JGNc6J1VvnO8Se/wiKuHLrTCtpq
1TGprhM1m6c6nFNkBm0HYECpu5Fj6j6LjB56OGiW5j0f6mk+/xgR/XbWzTOtwiFjcMoTOU/clSKX
9E9P+itjADtjsdt1TwbNciQ+ltxOMqdAohrYYmz4MTZZPMENiJq062T6P452eO+yKdql694pGPju
ZIJd49NwRzDL2p5A6Q0sQtLlQE11DTxyljuIk3Uh9zHqUsnjKunoaWvQ4TBDL/DGIQTZeeNZIZf4
DhhGshzuO+K7fBNE+7XDmuLMhnKyF2DNdo8cd7wWn4bk80+wJw0Ux2qoU2+p++YTsMuG6v/fVnsg
uUL9T5ywWsN5/jvKJUgINkqAI6goq2ZFkKpyfbIMBHDPUmGBxj1c5g9c0t6X9h+CQQuWaVK84Tqu
47iOrGxuUKlWxwlrDOuy72bz4WpEpXjVPwtf4q79JWYt3B4Ul6dIgUKMpIHuOgBmslDaKIpg5w/E
5PwiNcUlU5koOyKR8wjMw6GdQCzVfOJ9rArlqaIdR6lWUZnO1AditqQEWrOvx/cszmPtx6t905ME
lc2woy0tz8OCTiYA+FWjM48SZv+g/Ioadd2/z2SOI8JOsXxzYd76WmkUgJQN2X7ImQCuMCVeHPSZ
zWoxH7K7MJ8khs4Nk8koRY8d2sDdnbfCCi02da8KFDt+yVxTYwC36KfgVwk2IjGJ+9XPfHUP5Gpi
Eq3NSde0xqnyo3ccYz21Y1RWy/pkHR1dFCB/aghnEpgndHHE8uy5V89phsfg5++v1VbNG7/SeT5l
XsrpzhzgYyAC4rgeBWHH3oiwDqxcWZGyvb/8iNristZGMy949yzfNcVCyTbNFXaal9eG/uBtm7/G
tAIDkkxtjpUsHeR5ufBG7r22lo6PWjYFyn5SVOv1SheNzggmrrUhkeocUbi1jax049xlqKxalZ73
EP3HlxT1cVQpjZUdQh4lCWl9MnI5+X9lWtwxvatKir5TuMnbk6Q4uNdI6yeozk4pGr7K8QRAgVn8
PmCK5roVqbO4IkCP+GHMVFH4gW8SXGfPq4W8Ks6qIH8Id8AmQJaR/kESr0aXpqK+Gevm89wBhGfu
6wdTpo+FUDMsG/C2mmW/XbTA5G9kykuZFT4MJdiSW6CkoYKmciMckLE4dEyhU+Tli8AMEgK11iYR
LGZJtoKFdl1OiCjUbc4K9dUmKz/ldYVzULbcAgdlTQWbaBnCbJCTzFBNpOTg9wbCLtHzT2DHzto9
tVkDr22SQ9tq709mJNNd3NBedBYC+bReW3J7KsnDTMsbm+Rcdm+OHoaUeMdpevd8xb1kfOqM3Xbe
8NnHSUQ6CZiu8/fa45GuHMDzqgQAj4wuWhilZS6pmvcI4Y/8/kgLZeCaJbiS/lxLKY6O2Z3Paxd1
QgucUmEl6hBGGg7KSYQvY2JvWx2ks5OKiG3SWWhHXCYXS8sZIzmIpyLxRrWLuLkj2hMHlHZ/sB0u
nR0JZTyMcaZxEVjgKeNR9K/QjBjKBNmkd7rH82qtUULPqIVMYaiuau7mR2V4uBRjlwqPjBUPY6j8
fTOMzh0TaFbPvyUZGwPx2DI90pqxt81dUvkN1Z1PYJm7b8gMPg/n0XuylZDgMgiKKa8FZ3+9kirQ
jnzy9RHD2FkoMtxmj88xlgTPAbA+MEBSJ1VxFQU2AX9bTRwriertZ4xChavxr2VRcpUKOW2Kbncr
Lvvvz0XyCtGwSa0/CvD/fAXfYJ/wBva3rQovnmnpkdM+CoZRFhvQvIHDJ/T0EObPVr/0/0jRel/2
HNwa5hXlhzhvWLkHt1IUtgVA00KTxSiJUsRPcUBTGT+0b7Tp8pjq7NjtBpATmxiuy1XocA8FQLPw
D3XTdh2jeoWFTt/xsbi5YUF4PskTMkXdqF2FOLvMkn3NHQkJydPLN4GoTh4l+HSoqn8V+nMEjONp
BCsqAKplV6pft6JhADktFm0pSVp1QUgfvhXmnQe+G3My11q7g4lD1IWYjndgr0laAfUUXA0Lg3iB
SdaoXMwbFGvYQYCa4KBP714k137aqcs6aoW+Zwn0PGZd/lOXxX50KUwJZ1KevCcJQt/geZl9ozm/
isy0oIopJ5RcoK9kXls5LTbSfGC/D1cCEUaY73425TWOZqGZJA0zp+Bm3RzLnrIgGE94VR6RMHr+
kHKe7SVORXyRhiXqHAyIly2nhvcEQneudiLb+81P9Id9tlozRnfdQwRLq8c7s8nxEQmGTWhwRZ8B
+S9ETD4Ct99FbbSalQDM5SaUcwHl5cQ5kYXXX9YaCD2/Vy/QJa+z8niKQWfKXmIdbJTSsT2AGt6J
Fo+UxUsBrOXRwRAxxCvT8ZZNF++kglTH7V05Zb8j2IYRhL/8+Ulc6WxRDhId37EqO9vCVWHdezHg
DFqHFlVMRIg29w1SvA3FVMcGEojZyphtW7MIhVxgorVPuE6BuhrCCTI+xsDzXpiPcsbdPFTehc5t
YPAbMO6rpI9xISYUtiH3rOQhPUbgerrecL05lPP9PcgmKo8lnuCdZNnqK806j4xZoDqUMdksseMA
yz1YYA/KzGSZ94zhXyhbofpu7j0MSxFo3Tk6XC11lAhLcVSLdNSB3KRCKqpgZAybxN/ko70KvtzZ
TV9krL793Qvk3NohS/Z8eOSEnv/4wOXUA8QTUiW9sxjXgLtjMZbElL2zm+CFs2bqc9aHbkU9RgAr
gyIXBKJVwBt0TVUkKeIz4IuckbOpNDEms8ghLE8l0NnfDlKFwWQMI489SEySU1yu54LN1YHROLIP
bo9ISzFtd2iEZJlkLneEBWKIcQvdM80z/aeSKSXvp2ebAyykAZkbTFUMc0tQMt4cVuzKs/p7W7/o
TLefdGn67cW9ws6Hst/R8SF/JFPyS2+DAlYXfZ48XHd6nds3GmRyTb0Hxqw5+fGTYH/S7Mw9h5YW
l8YO1vGehh1qmDUKw6UbN4SZxteZ+ZpLtMQM0qw0kUVXpIKk3wKmaO/vL2kC7H9PRO3iz4EAra9L
o5UNtgmkZS2Hiky8hDTr/jY8ww433fO0i7OS2CywVGr9mk0O/qeNsUosz5BJcSMu/trkPXGd44YE
nvtasZPzXP8jUNI79jAzWFFkz+zHOQWmsg0dy4FcZ4ujQW7WFRBz/PHu0i8OUdIB3Aj67lKvy8ND
j3Fpgf5hfYeztjWUbRmo7n+O68Mnl1V5R2cQDdN7U2C9XoNngRMnW6HNX0i5UWOHlyuO40tkKGeP
Z4ohc5Mwml8wsXVLWThSzsvJbLNWywY5hIH32p0DJmIO7OBf16dKGGARmzb8Fnr2d8IEy2tFiSS3
fYNWoRkYwksASa+CSsDwRmg5ceegixGoF3zq5qxwuNlzBU9liX45bBh7Xb7DTrO37OJBmREYSEsH
OSpSt3HC6hhIQTvsvBxaZwD6tpGegIXxEQpzcQf36gl6Cnp1m+HJLIwHvd72zXmzJgqwCJCkWogf
tTjxFiRaPLOe7smJsUk9qr6qdUvhFeZA+ksvhAlRz/7gGmGN+/o8mbJ1NytvOsfGyZ6mbKWwahA5
oVkatOQ7RyOJPOMSLOYWo3GmDoXcSfAywuzP13TEFjcubqNtz6dQu5XQDzfs1xjLmy0hwotbqohA
wJUwX4QnOkdDPpyGhueD4v/aSQWfGijgiTfKVFazj36ti8CYLMAxaNFlQJGMszZ7RK0AsNNCT1X1
49m2ufELf/CLnabAd+85OQCEVgWrNdRc7Oq3quu0XmKC7OaUfaGkO1k7Wa6/TPurfzpkYqjiM12m
/CIcmQNzTeo9Px7WH+RzFtV+MHhELFt12/OMwadTBBPUkWsgMLz3f+n5PaHec9utZG+6D8XCLdZ6
JGcz8TqqrDOJpo2o5+CIJuhIfLFKv3crvVEoO7tPXOHzZRpNUsp7J6XzwVTIFst3Dc2SwtofN/hK
IwxVWNdmZTgXR8EVjlwHWnSDF+QWcYVrymtJ7q9uQmxPcRVQBMoykXbVMHxQgAlZIDI1W+YBK9t1
Bd+2HJFJdKM1jXvHNp8C3BaWXxQLbc19LCPZhkoW3y9ErC0MvzopL1oohjBf0dGfijs+m21DEBsY
yJmD59yUcomNjXsHQtphDyoWT1E+11SLEYnvyZntvP17gRzxx9iOplxryix55CpPPYNmrAAHHTH3
zxW3UbZNbSk1OL9UN361yL+NTNoMzE1ToKdpteCJ0wYHBVD19HQ6mqvS0uzEELJy/kxi3KCp/JAs
n4+9y/zpo3JOoKMpB7nAFXlDMhrB6Qcx5ZKH5WpGEtAXSOY/wHrZ1AlH/EdJArvtbdH+ZpENkZKC
vJ+NnYvx6tcv3RKfSfbZBXO4VDxck29lxm9YaEotHNJ7g8uofG0vlLb3eAgUAU+3VzORICZwgmAD
RwjVAvUKpP3bxXdCk3Krdg5UtquoF9V81VM1ej0czPacFg+FHeXLGtptIor//EhxXdAASo1UGHIz
HkD6aGWd/rHbZfmV6TKRuEX1YseWYvafXtuHnarAXeVT3OZW2JnPLUvSnDmMeuIaBe7iEJ9+VBAi
dj7srcAzdWS6V1EnwhdY95eoXEWN84xUj5WLm26L+ISNJo/pwHBCxH33pvcSLyW3vfQ86dDb9pSS
Wr+zDVBK3GyYSUm3xEnNNoXjy0poOIusuoHru+5uwEtjx2TqljERBs/xd/42CaDlEvnYc4+62T1u
4VIiKCCZ7dM5/u/rOSLQ2gn31hIA/j6T2sRdsjcoe9GtUio48L9mpGAKJ1kgZH62XnhEbLoMqvH2
BUpcT5evdkbObMsnryCKgE6fQwlPbh8GEqJqQtrNMRx3YanIV5S2wrFDhy6nyZ64NgKYdQ4qRJKU
xv+Zf85sdUGGz79nzMo+ZI84Lc3knUzcqFVFsjK5hZsms3ev/elh+27sM0mz9ji+whgsAyMTZLxL
pqGM9aDv4ACXLGX38sWzSm253/UA58K+UwSjj96lFXiqSw2IlrqzIk8O7BHP30ejQl8X7JFLYYbU
bV7GQuwgsjKBCKjbRXFx1Qz0007jDANKp43iLWWQ3OfH2yHDnWSmJh91Hezbe4Caqk/HDr20QUxW
/YbpXmE3/TLNtKOsdlL55v4jHaCalxs4VLtKvTjw7hSMWq8a78q5bv4gcVf5js9A8c2OUucyyYaa
GS/IaSr9CGUkGFso4hGDqO6LH7DKlCOafkldWSmlPcRpCHlh2AIzsBpgPnkU0BznpeNXFAeWfPZG
PxVA8f7HsrrL7N7Bl2G9ShPvM8b1bo7+Ovp+fiF2ma4atMhQn/HjUSNy6LZFhGEN8DjzNZNkqClE
J6jlcgUMCzei4K1fGjQT8Rd2nvPFPF1eF8/Wbw3LAMmx/IvrsU/cidWxYb+jTaWdzkA/sgHpZOXY
Jvobb6P8ChOItOn85BzpcpfK87c7e25a4JZDU42wVpnBABzkJroaNmWwnQpCigcYRDnl+H1Ti8jG
vknOikSZ5iAwqATzPjJNVlnjRFxf74qa5k8ywXEQpuxWvVCnMDqEHz6grOnQDK8H+t5zR0BHYq+1
DaoNs/oMn0hNUA9wN7I7ST4SyMSXvx1fJ800UEOHuRGd3umffJy/CGTvpu+Sri8qYHfbD/ym0BaF
qW5d6jXC7E8F1Yj2wM4n+wQZ7dNanQqfaUXQYG2glOjyCWB4qmfTojwuMblSY0VA3k5weu8WUkAi
zmS+RTthd+kGO5nxFGYpvmwnoOpIO6P0B4RMJrGHeCngLcwfKKM0ud99ftEBX/9RRB9Hg2xH+dPL
0ufRg6ThIXmC/3kxaCvBny3g2Xh2tMXhwM3eDOMATEMO+zwSeTt+1Gc1CDPKiE0yB0ia4zamtL6G
Mx0wkbIzJXI7t3SA2Qm0aozxcX6yJlj4epc5dm1RErKs/3XqPv9pEwjYwuHwiEkAZSkSLfgzZ3nu
L2m5mIn1LCisXn2je9Fvxe11EYUr9y9GBATmvFDm5YYTHr521hSooHemX4nYaeSRf+JBCt0iI4G8
YFjLQ06WN+ro3oY6Sdcsic2djeU5WC0NPJAf8DSPBSkeEOue5ctHaLtW/FrICyP3XIjZYcUnYada
xqCca0eMrwFSlJYldcZ5sn/rll+ZlOb494ny5gQ2qLRg9v0tOWUAWhN7LoaD8EI0OA1U5t4x5sQo
j+HzGnDu0HTu4m6g1GaQO3p+FcVmeHZInqwc8Tn2Wdo2x+/+lLXi/bYgMrmBvMJKGUBFls2URYuM
U2MdgGCXni6LBqDKQhn7pHni2WXAORSzncCevXJUX+CcSUjCCfIzaOERxP28NuogvhWxST3gDPBe
Eqh13iYCbC2imO67n62VOjo/515ivw92HOrHHyCer6DyCgRBPbVqPJYVZZ7W2vT52Z2OJmC0KE3r
+7t+Lr/rHlhnAxoXu4fiv/BzzrDZmke5BURCfdpYa+Ui3iszQ7Bk302l1YtblATVs96fA7sUJsDl
n1SSL6osGl6iG/WdvlSkVZiTRFQnz0+gNdD9AobQCy2Qi+qopBxhfA1qiR61zZwgjSEmLO1AHcgu
XY13T8Pux2VEkhxWpC+Or8UZrD2NQuh0Uv9M/eG5uNbJ0DGSlbh/+xtpb3W4Pi7K9LrxJaAneLDq
Hc0bGx0EKqjXgoc4gMp2WYj84z9zAye+Qyux0qBoVnBfwF7cZx2tDhrjJENUAPC4bjIbrSSZxgFc
yISwRHQwJWKnv8/D71p1HHuaE/uTRDxzF9eY0qOjpxmjQ5KvmX2UkVe495rQxIP1d2ARdgQKTIO4
qhMLDXFRWOla7iMZ1HIQaQvf5tOQ9sEDkF3j0ETZFJ80CvDwG/lewsWTzVlQmbgcl8tCDULLT+lb
/XQ1f/JbWX11Dpf0OPLu4RKh7UD7xX17SbYrBUDit091ZxoWwVUwcqQkzgPLOJlCm+tnIFSNEZ7p
qj/cLL07qfnnKeSUegIN8xprtSmYOiHNEQdb7sL2CryEqA8u4rPoRPDwev+Xd0mTdo8f3RcbBA/N
iLjcr6oRQW8CKTynLM72+KH3vg4BV8sXyQVHWRW7xL4O+Q26u1k0NLDMfM1Zc+LeVK0P+5IOcPaQ
PTmG2mpQkUn0NEab58d68Hhj0n9SnivkMnP3nSlDdrAybXHqFlNYAV2fxifisyYAIofATBU6Cz9k
5gIwB8E42HAiMmYIV1GugiLuR/kdWmgFvQhS6+6dhKYVH/NRVSSJjlytdeC4QnlmTE0nz/dzj2iW
ZSqY3YT5mqoFs/4+P295J5p5aMkTLZw37rAc84h0xOW4Flv+vG5sOG4H9KLfM8ozhkc/iWGuNeZn
SuMJwySXN+OoY0r4bmU7BKhzKuBfdQstJscBE1X5B1Y+HX8M8TxKSwB19gTRTEtAJAGEF0IkgTQY
tQUGRRxlHNd5Cl2V+8d+JD7hCUY64noWAnD29IAmMysZn1DtZckjvNfz5iUamdVJQ9rJJJx+zmlG
eEbotFlv7vhSZdFRy9S/YYc0/lbtCSmlm4PSLg+ACZbwzhD55oY7EoFHShHiHw5rJ2uoO+XDbXfs
Q6+sF6r36/m3fx4C9ewhQlb7hlrmPm1See4rJM0OzePnGA+XhzEwi/5mv1IwKb9ASk9vBAoJNvQr
WkL1j7JX39z4x3SwCAMIxZcsG8mWYTOXUStSAjMm7VhcBQfiPXzdx+xf3MBn8qf9RHKf0Fp91GkS
7O2trBksdDO/Z2Mze6bhBzuEpBlRQ8kjt08aQQ70vXLIQlxljA8zzx0UHhezj8Q7L09T9WPr3wxH
NXLgCNcYTFgzEPp/T/e6CmPvrXTIey4c4Svo5U5Mka22SmWzhKl0bpriG9p7knRN9zJCXHD3FVdg
7aHClLaKqGER4L81nfJguLoQXW69R5lgg8LpeMzI54NhChBR4+JDU96s9mRUt6eZBJyozv5A90M1
AObPzOHt2Gc1yO7Xfq+d/liRHB4qPWXl659xtCqIyEoBBGQXT4Mt5iUn2hL+WFGOvV3IEaRvaobs
R6nxieJ9wJwekD/XxfC8deZabT7dVec/UtPiBJeyVrnjMfN92JmUcHCCKzcZlbDTLJUgYf3IWXkq
1I3M7FshZUReVm2HkK2NvvRhKfRcyhUi+W6nmG5LHxbpy9CvGOo4Pd04tolXr0mGZuJncPhnkNVY
9t1Ist4JPjpYAgIEgVZHy0YC1xxTVJTZ/ae7FR+YB5iy+5QR4XLTfgPXtMirLdshL40McgnfrkWx
mw8cNzekZQrzzSRFpDfhauPzO1KzXmi2Xfe8PyjIK99x3riDCtHty5GUwOg4RYw4k3eQioVG71/0
/5xMi7/0LqL93wjHJuX7BisdDeDsxsJWaecfYtW+9vBKCxZWGAd2KzkOBUHrkc8gLbenS7J8bZbA
h9sk1BLRGvZxbiINErHIivpBBYEPYjBdnWAyolj+NuF2rg/6txI8yrOgd10vp39NbpI1CEcwxJym
nptYjuax5a3xIvmG4eao+0slB9GlpjV0MDcGWgSF1DDnmyNF2KL70zMxO3GL4RwQzfxyms25dT7g
UhbCzUFvY6PV8NLUz+54VTaENQX2vOIrjYdt1IqeQMq5NkqWcv6pFz1H1eQSDbvsGuXzc8CXNzLR
LqWSV7l+YxO5NKOYcNYYrqEeDsqJ4+GJwKW6SZkz9Oqa8IvOYSfE2TYiXMA0NKSm9GZ8ZtCTyfpj
4q6RGS0oBvl8PIiyUoCqnJkcJP2oQoJjWef46duopcIM9XR9j2/+MrcyTEiSAG0tW19SG+3SBrbO
uSAFnJxrbkLzaMcrZb5N02Gw/roEzcRKRPxPQz8TuM4ChqQd3xE+PmgJYEgXT6dLDEOMdZk4vZPJ
o9nEeDGJb0k98lZSo5koI0ISj6ghnPaYlwcfLGFLe4rQpmFYvw4MvAwELMTtNW+lW8wl227sdnBE
1/dYDeAGdgwpm67H2mpj5qqEAvQu6F7x9C9GeptR5HtCH2TgK+XF8T1zNrUtY/zopGihafDNGAiQ
tR2fIUAnAgJbTeg+Ri5PI1pqs8wE8tz+HORNdz0cbQ+4cz5ron+Zc6F+muq9xJtsBiRioL3hOD/S
6MfFGbdTHognffg5xBphwO8kLdhTozUSRv5JO53DqrEvNxfm6XjM06nGOzZ4HNDz21t4wmjFuXz+
RYTfTDCjPJzseDyU05VgG+sAO5D5joK/kvQBXPWsO6fFI6q25Ax3w47JMqMOrhgBxa+HQmBeTUo5
fcucDk0tJL8wcWmpSdfZLEe1BmCOsvX8ytPw7tu/onGBpLhqKpQ36nuhRKgV1/tkZLscphdD78CI
5enzfxOS2L2NTmpMvD/oHiFl7NpHWIpeVHt0UW12sUZ15fmovAD3JPEhQNrJkBnzwZWgC/vg7eu/
YkWnmn9+X1w6lvC7JiNsXSfVGFQb7DhsjdmJS/9rfYT1+48G1WZCI0XIRdiX+5eZzJMTWGmVnZq+
ZxzZf0d5sN+rXsll2YreScmg1TvrR/g555MML7dH7AQwEssSkUa6EYNW6mKUrGBBIWcfJzJgLdV+
lQdRLGtEmtsLkYULM2azq11aM9N7Fvf0DQkj0gcnL9zp/jWaNE7ZcPPW4HSv9OgTP0SSTo5JUkgS
oXUSTGPPQLbZJinjJyZeVNUTpcscGcl/v9kq3spGJ/BlvXpZGRN4SDPIgkPtZj/UZ4CE+wdotRwL
sGtfzZmumDBbZtquin6wz150Fxd4E9m8KEH4/oJAoHq+qN1OGhkoMgT7exiLVa37nSaPFTdaaRIN
v9uJ4ERcKfulXu2N2da4HQtEr8NDWkM9eqgAnSaBFIoPp6kGoSVBl2rQGurDC3MIQ7eFNW39FLCW
LoEOavSRJPzW3nHdxBc+6AK7mTXA/D/xoTKUG04EOoGmZeX7UPtQHzRhc2h/glBMbczEX84oSF5p
sz3fsZn14CNuN35Kfi/RDlNH7QzWNW79+bd7nIt8x9GggLOiinLH2F9neFa9I8ZEJvnV8Lp3IIBj
oIkNzPD7kMjB1+2tiFB2dWgPMD4f/lhQvmZxcBwGO5rjCXYs6fOXc6LtyfoFjV7iD3sCSv0LCDhe
y0JiyOPVOPEGlMmhVr2tFhc0mY8Q3vxeppMZSr91xU0x7CACk57YLVNo6PKXBuH2Rx5JrG4bjdLJ
fZd+hm9VDq59nEUGPq8FZWLZHl/1buvV/jEGVNWerDnqyux8MN6NChUQJrT9x0YHL5SCYlAMiZq8
3eKKbJEfgPxuaL/oNFzThGFiSoi3oPDDMuQnvDz0GEwkJA/rS7RnAzIZHM8GXaU1CrHeAwivyMZH
UG1U0cws6JgeJFEgItbkVVw7OpPqJzQwFo2uVgQdSBiXIiCxKZUqss6e0EqAFDS9Rr5dSoP+LEtg
TELj4eNMhIGax0bE6LJdGFs3x8HWkkJVfJHNKCtO3iTyCzA8hWBSf4Qq9oOJLOg78+lqF5aMpcm7
EK+DZ1uf+kG4gWzkq5mHUMFVdILaBJo7CP5+R4tHQ1PfkiF/ouVjpCtgZJ5e+0lxCx6Iml1nAQ69
IAZnaPSk05Xr8KOG5pK7Y++RJ4eZKNPey++ygoecuouCHw8OVHyFEGM4GVvc6pSFmkxvCpq0fUL7
tTkuh5024ZXVRGDBThQq7bOt6fAA6lgnglE5TnSP41iXXbCkky48A6BR4vOBaGTWqqGeF7hs1R6q
a+thw1PGVISndJT4bYQdH2MLcMskSThYWX2woub+tUM3QssYNHJWErP0YliCzeR1x6/b17uzFNx4
+wtwZC5m9kZ6YTM9Nh2nNE5E0xmSdSmWLNXtELY2e+VFdobt2nKB767CuRO2XWHfGT9Q0Tmz3OeH
x6SNSOiftF16gBN6yxpe5kRAeXRE9KpJThLD9Qe7majciLtLonCFrAByLig3QZjjfln8N5gEpre0
S4sOjod0BSOyYdUD5BbCa+9YtdZ+BIP7XORb376d3IhSB1qqmWVg7jeHrsX8WnaW8xE6XrULfeTB
sJFSHOmyxHOorn84I2HceHKVyMTzCNzGWWQryoE7NxmjqM2o6posN/1Hia5nglczZgv0ytiBrUx7
X8gXEKTBbi1jv58ovAP4DdWyDv+a1G1KrDMbrE9Qn9NRvjSPIz1UrSIkDTkhbSG6kz3yjz86ErSc
UBCi4hYQiSjXuEb2vFatVs/zU81YRTAQRHXQChP3M+C/bPsGpwRRFZSrdbXDs04PltVYZPpcDxl0
bzhieyJXH3oblgeH9IUDV7jS4e1KVUcY2EbwtXC3raP/MoYt5wux8IRZCiBHSLRzqbFxevyKgjKI
81t6snI6rSUAplBQDVPJl9LOGePC2kjYEexf7ISfbkD9vNqZtSF1ra0BD6DTT73kK+ZZVGXZEteH
HcCX2XXhxx9uEzjqH4nTr7TFKdxldhX37Gyl4XcIxnio5GXaZG+0VxXBTIM/elvuqIZBjF3ygKAL
TIg/xMc75+UafeqM4BCYYXM2Mg7Rdr3b+VbNLxKi51KS1qmjJANO+UK95kNPVbn7UPclYscCKmuw
nlZrT2NyxelTRjiBOlhYfDzEKzDiZKZaP0hkwfUZ/ESUhZRQbTrXpDLYwOPN7VyVjzO4xJQI7/Df
yBxT8is+ElZIIRhGxkJW8bNrdkIxNesGQ3tW3y52F/qGH9COYnZp6yZpXeLnooVMMfBgnuZcFYVv
l+QCQuUk0wImv2xB8JhPfwoZkaS5FkxW/UfUbe5xStJnAWtFz1JT3PZqtQa/3DVVQNIJXaJMMoeB
AMG+lhif6ax70QPX3ly/NjTI9f5waH8Ahs4g8H6MEwIIDDWfI6icOwNI7L8I2Q1q9a3odqjW2Asy
1laf7YyRIlwzcoK4Umw/KCVmNVFoO9iIVuYDJjBnockaD17PDVY4L2vEWFn3UHLZpRaDeTli8sxr
R3nMbSpUgqvq5ieeo7aEhd5K7Mx1OCNfirX7yVzYUjOE2kIK9IeUK9mUbCq/dNW3H2T34ta/mHj1
mu0a3RxJ5+vyydpcho9X1wlcLUL4Z9KLWNKqTskkAIzk6p8VqxlJCqMKKYQ4ZPDtzR06DivUyJ7n
6d0QAP2kB9XT4hsGN/0cWEQdSNc3aTr46FnjfcDlg7sE8/XsOOVj70DB6/jC9dUbygQ7nN2MUVWX
7lNnvUCMYJ7fQZhE+wLPqnWaguD6GVnP4gWStNsBj/k5LeLewsn0hi22z3ArtwauRpRhhJqB8WUk
5uc17eaIPLTIHkqx3Ci0HvwPP95kTt/XO3Tpx6QY1oS+e/r/Kp7H8qx0BgMzZ79wdRGekhpi1Pqp
K+GzwlrQp+rpHrF9S8RlsXoxVIaX5c4C+FDXW++vdyOLA0i0qMXY2nh3imhF72j7G3eCP4kVsnsM
Eiegex/6gmrPkuqivDQsNLNN6SW9qGM/J+y/DWDj60FtD/K85NybOtdx+kxUjAxAGsHxaD2wKD7Q
moYxnPVQSPfYfWo71KnBgX6nlcY+nbEQcT0fNPi4ymeNGlkarPKUa3+YvgTQ/AFaJOmlQWTJ/jL5
DOD+s7M725EnCCeFvGbhvJmlbnrJzAW0r7icoyxkfIo4iPlxctS3W4cAt/tlrjU5NwHOIhJMeO+x
+hJppj0jQhOsn7vz64kyGMzrGJ2vbSP0Rr4K/IpWK7qpCaZvn92+IZ5+51uERNR/3gzclmTms9ap
PsHTf0NjmgTga1/bcohk+KwM4C5nuF6sWZZ78AK5AYUwI25Zi2KZ9aW+VEvsQKG7vIX/+O74XMLo
51QuQIdDoLSbv9z7yTaOLDPs+9lq+9sSDY71LvY2UszXog1cmYGjnf7VZ9df0fM6jlleYomyv6b0
jcXxmay3EA81xUCRFh63EX1GBI0R3L/kW3z0ZEc7KxPM2gaj8uyDZlUu7Kr4r/RtnGAPJVzsTb3j
3WB06kZSUIEMgegjyUv7S2RFd9upUclpl5gbpJf0JQP8rz28DzQthDP4D417CSaetndsgdblT6R8
+tfXeEETsnFEvXDxzTE000oR0raZjKDHulWxwzgSXM3dguiHIQlPma6ZCurkmPAzqg6k/iuGHa+X
6IHTmpyRaVk5oVFI2MhOhprjIRc3Jr1TcL5o+Ek4BfmVfdUh2ZKRYGFuje4b93j1b1Rj8aOh3Fpt
Y2mOCYz/6j6AgBjTTy7SYmS397apGspGRoX9t7NKgAySAOYoNJcGl3F75Z7s7aFetAOP9IbAuh6h
YLaVPU6TgHz0kcF0HazlsTeeneypFdyNwFSxnoH9XAw5CUDWJ42yqI6+pXqQImh3NNQnIr8rIVI7
NeysMS1Ssr276jd9B71UQyZS1eZtV1cO2Zs/MQLR3We7ILW3twKpD1hG13S4lVqN+2TD2YU5BiLp
k/aaRLIhdZYqfTwDCPJgHIj24pNZHiQtBwZsqwV++QQnPPeAd6PRIjLpxYXQqyMasAlyUcE83bwE
F136fX46wKVzv3sas26yjgi4RVyuAPz632TmOU2CfqwKNgRRNgWM7sLTMaIPH/PohzOTzF+zREGz
kc/8c2nzM68IUgUqhiAkkQ+/X1zV2p29zxDf29Oyf7zx/vBugFM3IuEysFAxe+3gQ9obX3F2zAjc
Wz7QstnYY1hzRJ/BebhRiQPdEjEf81QFIv4AkI3KkIB/kRjhKXbvhXMiacwKeg9mBtLWLU339N9j
pqJJjzNQ6YbHGCI0WEBsRVpbcJM1j7LQW///lZf5l76vfJyHgW6w9mAV8T2t1M7MnRIxsNAFwGWR
PTKbRIarBOvLYwV9KPe8Afp4Tq6N88B42eKJwN2jQJydo4BhKwHeEUfQvhI3E8QYBCJBaI4d/3H4
OEVHLh9C7lB+HcbwAXTk+Q40h+0+oTLcf2XG3hGtmCzHiemJ7KLAVZHAi6UIr0ijmCgRlvKlbX8q
NMqJOhmhafrapgr50mO8ZGyM3cFHW5RlKeeiAZAuQ4v+7txXWnuSaWVMI6tx0fw+5KvgWpzbn/2m
V7TPW+Sfqn3dwtsnCNnEcR9qz4M+wo7khBzZzlucoXM+ao5BpMYK8IKrFTyVNCZkofMbjv4hyLw9
Wwi9JFQQEUuqluaxDqNkFoR0ZrnCMYLFRZg9u0s9NBo7ql1rEtN76/oa05R1lNMUs/D2cG3jUHKb
Jp10+bG1gTrdxAwPJAq+ontOxDVEHzjDrpRJPykUa7kBMEq38gE9ZOfaYWaL6/kmrHunKFzzhV5M
mOcCic4yJ+ut8eRlhvFFo2+PlBiiUmFVSwPXZsHqGbU+/3+BvYOvEaQU+p5mIti20XFXLXc2qMmP
v8UXmYbgXhCctYHFQL5pgsCBxlvX6sr+b4TWIAlIrdXySsmXM9pxr9d6sWQftHvhCIBCbWCviwgc
XMIIkl26pPaxRFr9p1l7KbKmjA5HK0g3FxFOJIsJGkFemEvqyKOWs7ZCCDCVEKzwlQ1BqZayqSUk
yTpNv0b93l+K4W0kDRBhCZk7xFgfD7xUV8Vufi7/L3FPZ5R+ulTeUS3ikXclyGsWYcx5vWieFpzR
KuYPFyZOsbXdD3n40P711Gw/7W41C4Zl+5iSkDHSrGCS4ZbQbDkQh0pynrjr5mcqMw5x148ftB12
Dl1dIco0kcq/99wGBnXfs1OThpGCt4dWTWdgXUqO93UeBK0t9crmTYDjh20miPoABuBRJbpSpKxU
+2vBXWQKAF2RM2ZPSJZ6FKPaDfEf7wNCYYvdhgl+phtdck99+5uiu1h341NomkqrF08tNYY2xZMF
p2qNE0H/WrgRwEC1Lz4hFj8y2v8ldTQMJo4SOL4qswr18UxGGd0zfdJCliPsPTXWZiDaZjUd1JWl
j+72R6E1yIj4yW+kuCojU94m1TXk6+Rtv76twsKbh8DkQb4gSC1UJxLMeYoWdITYnngLn9oQCgUz
cUsediKgLCWMyolgwNsIFEF+ZG7e3X5Gij/Wx8j8KexzW0lkmcCKQ4GY4sxBKUeLdNSZsB00JZ6r
h6ltVoIhV+nQ/UDRsijJFB/Ou4XYMolKA1UR9QRS3SpdUpywmVgDE9Pm4C3PGFPOKkuwxhWnWNnQ
rIqvJwBCigACr4y6hl+G4WHsVRNUXpXejF6gzPfCOWM0MpSaZRZNPRGO3y/xogGvZXXdRgDwBEEM
mwUV2Hh+q8p0ki8DNwk4rwEZEltTMl7DkyPyyoZryhAcilj2yJAt0rZ3+Y38fwAQHcOXW0QIANTz
0ZSmxyIzIIvjE7mYX2JxRzekTn+SNUrrN9wDwpwAat3GIOhaAyKvh5l0G8gj/CD5t9CnfiEZZlxU
ZX9tYJKGxPiCd05NfYPpKNxbEgGeYOapH5/RGPKSidZD8F+NcNSy911JavFy6cqTPr1umw5gphsj
YzV90SpJSsLp6FFZ6qtG0j/F7Jh/YjvGsvMYBBfn6aeyDd+5NRkHCs3A6klMi1GAXZBMfXxVJ2Lt
wD7dMBG4MTlevuzcY+8iemhwmWaPHLcCx/lFU+nImLs4j6aosmnOeU/ohxFc4kp+pcovN54qfwOo
rJCIPiJbXIJaVXaY7pv+wGXu5C9KVZZCxceCw7IF+KMSLzfm8RGfoinD/Rd33gcz/LBUauVS8f+W
budySK90hJPqlV6PohMIYY5by6tSgF4z6w9fsLXiapkuiCUBSp/aRKZArP/LvBqCQohD4CDIvf3A
13IMJJkpiSRDBkNs+ps4ZIONQoCMAo8/pLxN/9iZVSJ8aWmO/A8hEycl4G68zl0iletYie2ee1gs
AvzSy3v9vcNGycVJ/GochEWT87Y60IcMGu/rtOKQVPSqxn6sbqnTzGLe6EMA7S7yePBBFrjcFWfh
filw1J0lZzV5iumrAZ3721EsMyvBi9vKN81v4T4732wLi2hXZ4qR/50zkJ5+aKaYKeChFMhi7btA
1AuMOCh9/72r6aHDBsixEMuzft0L41A4rWZITfa+29bdpfw+NgAmDMq8lfUJmxBGCo5g8+wGQQMg
yeCn0gpLB7GGxy08chEk4Pf0u+ETf93WFfrUBDMHjwWzzU3E/blFzEuyRjq8JHPEiObk3DBv2NZV
KeXcOiJHx5bj1hS4b6iADu6NnIIFsHLe3VyFelO7AoZXJ96fpPU58P2hwrzac1Ni9HNim8kbpfxB
5/SKqOJGWm2YaCRHBIF4UvnLJol9wBbIUu0r1kh2gHol5apZt28JXTdbMjIl9CsbHMzVa7hrpZkD
1OrqEAFjeyz8Lw3+/Y18tsHoHjWaW8EsRTfgdO//gKTGvYBzs9Hu+CpKpq4thOiaOcIrduxq9DvO
3aJ03IgqqW9TV2p3U/bjqA+z6rXdpTqtjM9YhLTcnYeLi8awuPzNBgW7HQt3L+ze9C0iUHSN4D6t
4hhPct4cWB6YvvsGXSfhcD45oGPj3rQlgjAe9w6IfDy2qVn3q9hHiO1kvTPdSY/RDOveRtEFuvbB
q0PqLn8hDp8QhYWGA+G8JPVu0K+IReTC0UZNhSZv8qjixvIPfnghnPSRoaxHzOgWOrc8rRHtOv1q
kRBs9UXMN/QL9X6Y1r8B7wRPGDmSb9NRrPN5Y1gL3EstLXy5xRDJkUEIst40bDgO2zCXxbDTEJxh
B0MqWcjdYxhPjaLkiInHNEFxC4M1pZ0LbWy/0wFsSgDWH3nhrKek1nj8ss5JbcC7oRxGPs2kh9oF
IEhzXFC1J46yCkJKd6J0bu6FwImI4S+rLqwPnj1K32gpvDlXyZoF20U8VFFi3ZtSsP7NdNVLBpWz
gI2L7LQJR+tVYYSfkWsqqpIeZRHGVI/HHAZd/+aQVBAI43I8HuyZ7pDNEg2gmYu42sas6NQRQnHE
Oqdy3Ft4WSarnPHqoC9Ruw+J9KrfmVpYLoAJWkQJ7voSxPT6WL4Fujr3LDtn+m2HIKB8JOxPllzQ
vL8dPr94SOGn8/I4xOUukX68rqpdsmZ2YUBTtz/gbwmh5wk3dzqg2ILFBMDaqXP4Lo03dBZD7uGX
jGAGa0XocoaXNrlZfR2FhQWbqBRx+qdT814yhh6ZApPmubWgWQIiTZ6lOf1risRNxxnSioM4aHLZ
kncJ0WAzc0gLT8RytLxJsp92OOIwh7V/TKHMTLz2h/dThE/4vwUySAGcuN5I88X6XCbDTgqnscVr
KJ6iao1RdrAB8jaIJrRl4SL3AM9aX7zWydGNrYxm1nMhqXT6kGXZi0SD8C2eem9kOjXRbpIkp8jA
+zBhS/h7TLw7FopzgekV7BXBLeP+rRuWXgCFaL4kQgUWrtzXBJYzvt+SGBdLsWmj5Vz0KE/TvubK
BH90OLmizY6Y+s1RavFnoBOd4duzr6YWEPBq2MzeVquozhY96+kwybEzjiSpDYCaaNXGS81yjiV/
raBaW2PY2rLfidZ1EUPremGWvF+zhTpnYzoYu5oiGrHD65+kPhVWwFQ1WMNsacMD4xckQ9ZWspmY
3cql/05Mof11KrZ67YyEF5t6ux9xuyhHpVv3Tg1B8FPsKu4ycXxvvTYZPI2IfX7Sj32MHVh1nFGm
5YAPjCOOm9rKIGehntSGhtcgUh2DFlyfWa2DseHPbrbrxyKoAmwXiGhHFM5XvDqnBTUt0HJ20iUo
AOpANxICzJyDCQMWbgL74f3wYERSYg/qfSDMZ6Tc6OYH70hqkG+MKPz6q1dUCvwixQLQyfNh2drR
tfDpRaK+jVW6AwG62pk2LNOYwHMy5M2nW53g/IxodG04kvGEWOhyudCXb0qU+z3heZI4BYrc9K2K
ZQK2iW/sJCnA/kBUTyf2U7WpJulmSZ+oS9yacjQ+6engMDnqovYkrvGfk+rZzD1P4xvY1Qi8uUsB
QjKcoTTkSPZq7VBWTfjhcOg5scq9Q0ONluI2sZxOVlSi1w5A+dArqU+YX8dGADcLp8CsiD9eqRA3
pfi3WdSpqSCQ92eac629VCRvePFV5oMZD+rGjqiYYNnGNDJm2dv8ts+F1wpWgYOq0j3HUZe4zoNv
DKhp95RnOAfifTz/rzvDOYfw/GZpupogtcVC+dqTkEFqVySETLQkigCTdMG5f1qP/jQcNT1ogYh2
GEXG4eC5UHNnfjVSbnv9PJQ2AY0JNVw1Zo+SGpUPSe8JaxzGH36DwoTBBKBOD8cadvBXil8LteEf
lYzgaPcM6GhF74ya2PYv1yiFD6A61fxApyuHwusxVsKY0tIJEC/SUdohCf7DrahpjK15cjMqvVGj
skcfr7Af2LDBaKtQhrXDzd0RQ1OsPHNbP2InAYSX0eRQhBm7QFx4lWPHB/FEeSbjae3U/sBy8rUD
7i1/JEJwzIWuKc65h3FgcmrvUW78wVPqq4voWjOnk3OROgHNQWFqtSv8j3b6oftp0B5yVqVGwWqL
ORYhYuEsprfx3FHNKqap7pHssh+EPMcNIdpFLjiXhMGfZAFafnIBkrjPGilKLFaVI0q63n1lBEqK
eURFOSUWtWCGZoUU4isUGEYT6T5ef5CUMRyPc/G7xmeGAwzhdFXH+iZRkbKYn0i9HT1GqvW6coEh
MNvfO8BoMu02q1jHgywvOo2OVxyve3FX5PO76JYuKrEfo+lIwu4Zum0hTYuBTjefzvUY6LhYxhCz
cb0HH71llsR9E03DfAPeCvxQbg8xJAB4Jojpzrp7mUCnAzmFbsO7YDrYQfLONNc7zTjKg6jff04b
ht4lc11pB4DawdFJAjZimDqcTdHAtRZ17gS/SxZZgSyXsJazomWzzqcqWdNHMA/A1oI8o4zo4uW1
Bkghk11yGPDyhWrcSmHST41QgTK2YE+1w48TGM8PvtJPq+dqutEkSSMcG2Bo/9NS4d7A/xYXduSC
5LBlC9lAqi0XaU2YRyX9TuOMLIkTldW8v2iVNUp3pC2rAlMvYyz8FyVK1dpcBTzE6CvD+mO+91BL
zNVFGxdGrFbvWuyT6UxYbi64p87qS5w8HAF3NG1V6QgLnrXwOUNPYFeGks5MAKeJhU5KwdjGOnhI
nn5wOUUpESRWGXOVkc3kanjl3RigWf1pXbswruM4Aa7jaxpflwhfbau0feGvTR6kE4zdYZlNgRAp
u81vd1CMXnnV+hPj2ahwpFMvDi8Ur6jCrNYTIhg9+szYG9FUyMnmqbDAKm/7UH0K5mW7+tn60jNa
w5Wkv+jPVtkfJTZ/B48JxHa3+X9KQW8Kgs2MKONrFzGKgXyCoJOZ0lmndrFwI4vnmkHQsEVlsuaH
FpaE10iDqTnXCcY2a4sOYEK2D0gplKk3z1W58mVJHVyVDb/DSfuBZqbkMAsyDNX694SZT8I0QHwX
szjDst2Yia5idSRE18PNHsk9rUt0TizlZLRfRwzJ+RLpG2y4CnV2E/BxxsLsIeji+sf8Xqx5aZ+Y
jlKKdC+CYpMzkgXDLs8Lde55UlcM8dKO00WAMirV4PQXYX2/tQP1+xlsvyYcL33L64tAVV+8fFm7
kehOrhApOhZ9ZXVkW1YW9Bi25kPA11+Zz40yj531qvljQYwkZCAzi6YxsLRwmcJE/o3OdhmyBMpo
cTZzSOCnw7/m14gdLAvv37UVQPCFRffM8IcQ+uPO7rLGxiJ0jYkVWZvJw30z+M4mzQsBW2sG+uUm
CfMtJ+N/8JpFGi/27M/gQeqtYL4ZXhAeowI7QFGYr+SJ9RgLAXkeIuqc+yI1KBrzI+IUfP9UQT3H
2p3NZyA0dsiGHnqs07y5vSvTxZOwFqcB150HBVc7QSU5YFdwKBNr4o3BcTowzky38n/nWN9QL59k
/xyJl7hPfnHp6JskzHlL8edkAkBHrxexWe7u6zcq0clDKbSvUBpo4MoN71P1FHw7GIj2L1GKOioV
KRmtWfz/71yjHJeWQYnQKJ2MPyiS+LscfVEjiDYnB/MgjUMvJSKG0S+tYpExGrBl/nOzFMocnjrb
NmO1VC6Ti1Kfn6RmAiwpzpWrz4nnNgPnJlrf67Bvm5A4+R12Z1FLdVqgjPozc1Lw4X6VtIthg4sS
q7cxgm4hdxp/pOpdtaMLc+TLG8wY/Tck6pWL/9jqEKi5lECIwMSceV172+OFQdz9p1/TjwYAKqdh
/xwkdGbb3gFRLhO1CzQRzjn4MIJKGbxXKVxpn1v+nhlqim7VVKvf/2zi5Octgn2c5+K4EyARH/90
HOpTiJGirEqCX3/lF3IZZRHmc1G6WqdEryREDTCcCPdE4pOJJzPTnKzYt/Rw5s1aDnxfcc5KKmrg
ZwXali/1fuqaFt6c88rdidg9cTgN3l78XEwpr+foqqmFFIaRUwaFd9rffXyDz8q7DEYcuYAkYrOH
i9d7SWjHVJ1JUDwB1RmBM69a4WaP8Q0UDmP//WlWgwwmzUIVYyDAknpOZw7rKRKagLX35hkPB+gW
l9HxBpfQw4VPZCyjBC6uxGrJIdJVv7L6wmDrd4S3BFGRSevPKGd7U1QwICz493QWvM/xEkjExUiu
uu7M9rBpfvwR+fUABVkf7o3ZLmhvoLWsZPOSbXtfC5fren9K5ROeC2PFgUDA+uMIwUKuvFW+oFca
vUpHgFtqr263+9Y0KJ2SPglAlFayrfBzD4v0dss4sCrkfrj5P07/fwVGC5pf/CTao7i0n6ywl+8o
xPVERH0O61A+nVrxGhaXn2guEelrl1z29Z/eVbRqLbSxzutVgfMABG1E3bUrpSoLGWsjkQTOw2vd
D1/mms0igzlHr2UBtI7DUU9nVL53o3/1CUD8gQa0oJOKO/Y1tnH2kwHmmhAuMq1gJnw3qyPGvE4v
dG9A2CQ+kkLJ5BKsiCXEb4GHmHHXv5ET8v+BmLO+4W8Hc/XPLDduyrHxHTk8JNJxYSGA9OPKw18D
bgaq++21AwkJxS0BU2jVdhGauGIF2FpYwhgCxQbvRuJB2FeSfQA0ml508EsToIV6rK1WXZDE43tY
6OzDtokHuntIDvTkjyd8Sz9JA0Sh6pmXViaFlb2auHUd79BqoWA8FnLbewPOsL6BGYtVozKKwegq
ui96Xp2eX3mJztqvsNIMrpOhm2IXpTrkHamUUDqUmov3YdoPv6as7CBO8BG1xzwL2AAoRC/wV1HK
n+WjNBXqftFQxYlsin7oDbueqaFTVHvYHmcqmFtoxX3++bo1pRsmWS3mYklGXLWtdXkEs/4Mfw8H
A1n3wmOuPhxXQ4ttyLduUyv+0QjynxWxzbi4R54Z/tZblThthD/q9jI42uDsA37t+A3cyiBsBdX2
bVEYvMFx6+trn4EiVF4P09B8KW6HKkZ2/oFzsD5TUZFfgoaTSkx1Cid9X/MNYAEkyEa9kuE3BAPp
2LquaIOj/SRY//LQBVC1mlYbfqOYJYMuSC84ZfKveoQOZf7TOtBt6/qZCe28XB1MAwcgFkEXv18+
wAHY4TWoGKLrswjfmXod2ptjo5BO+JxSnyD1NDPrZzFhYwEH5g9Z7vBC2c+3iVu6P0SDSKkhn0u7
/nXePVEQq/3x7p1IVBciNTDf+CwUX9FICRxjG+4TxDDK/jRdNIM0R/c3OMLZUXb1jCorAR+KjOiJ
XphOUXZ4Y633umyTlYFsXu1d91sfhdvBFRLzPCVv7axya0W6BURHhtO28ttyE+RqUq4fRTb5o2Bs
gRCn1HbrwN+6PlHcULfjvlgdF0LXhQGIyvdmcAFgyq0cy9ANxxFQ6m45oEFeJDGEMYvdE9uEG4kj
qgbCvQOx3K+844ZsE2ewLCGKs8UeV/f+gieb38CJ3lYH/0G3v7beIpJfZMDlnnGi472FqxVIt1fX
ekO6l2eV/vbtO8yfSvAUP0aY/wiyov9lKrlVCTF3psytLWp95Ef5bJoQWk4zlekqVZVX7NhOrGJY
sT9hUOMrmbG/3btpcdiGW5WlzgWNHwSkogPyPKwCbr1XnaIEzRUSp9KNTKiHg9hg9qVoaHckNqD2
AJPG1XF4p4nHY5bSpnGPgcd+dBeOBTsfCc0o8YPQ8z/VCXX+TSHd8NzVGswkIF/ITxQLRYMgLlnn
Ah9GtmXpcMKq1WoLZhrobWNX6NNf6Sf9K71DsSX+BDd3Aq5DyKLiDUzGb3DVdY33PLnt/Jau0zg+
gpSTJAqEVhOMnXP5+h93+TFaKv7KoAufCqrglhlpsRFaMBnEVgkhtZhhH74tyRmRAzF1V1U5Rsfh
wAfL3ZpVRHqdrU9Ri6ruEn5YO+WaS3ezCXGqUiZh2MSzu7PaBqF1mveaHS00LkLREvc8AtqxOb2Q
hAPXiN9Cl9ZuP8mZLzQdMAj7vAkNGTEtg11r6tViYEa+Tf958CihdBAGR1R2gMgMgDEQKXx7phYf
sIcQXj3YwR63hzcso2oTnk//EVUTJCQwCQXqAgbt8Em4011J1J13uadWOtTimWPgjZpiaSdbfu3H
tst9kkbojRjl/xci7kD3Kw/Ls0h/QGwaBrPj8vy+MP/4xGkp5qOAjn1YkuVrY7tzjIbpPjgdbb9y
HWfVGHkK4qqyhfcRQpY963xAAEjdVv2UGmrZJTHwjVsltCG/Y3qseWPuzjh4ngSok+nxoYjcumWK
e0uOHpOpX6dnW9N8rQHAoyqWKDVjKv+zxWPxn8c8XoTnQ1RcsUGcHHoJrIRn4v6pWTIZr6RQuNWP
Kk+z/bCuio7ufeq10LO2KIqBXpsNJuksq3l7V5E1BO19hXfQxYCDC1PENRmDpDSI16Cizytel5Nx
u5x9dmZ/kZQk/Gb5v0KmTu+1jZb21rk6W3s+6/T2wspRbzEJKfjsB+3xLdxLdLMJ3v6Swq8zP3cO
7rNQKxpD6KSZh6+SNa2KzOm5gRGRK2ic2B68sR1fb4l9y/YCTCk70MD9qjUdnx9BY/abI4EYWy8X
DODq0gCroJZA/7WizfV/aK7ELn8BqU62g6JCNYLW/3w/t8MfdhUCAdukIZ8IKYih4CUWz6clwJu3
FF/yMr+x3DxFgcO5LsPx25BNW808ENISxGAeQY63lcxg6UcrjS/Z4FD3F3nZCp1r4WaOFg2+lrZg
8xy3OlGCsiucPsA+26V5cpYe+tMHmkU0VKW1noE24pKtThAba4M6Y6ZrLIc7jq1qI00vofQDK7V1
rM/o2zEP/csG/RSoAoMav1ZVITWj48lF7Wfk5ZiFpb+nwJdyGOdPE8C20jsUc4rpXRwbXMK/zgl6
QGSXPhJKgs2yGZj9vh9wDxY8qlawYr2naMnBA0yS0g0bF7AaNXoDcRbtYbgCpwfXjVJRRPjGMtR5
W9bdTQav8bF+pfeXhugGMNiRs+SKjjKTFLZ66UkG9dg5eplDf1d4mEP+7b5+9LtYaZlLdRNqRGTv
qcw6CUh22YG+fZ7dgnXwf/iQIg8d4u4L5ixlqk719iG5B11b07NA6dKW0JGoir2NP6o3qCVHznOY
Qy0ZVpSmMrvycqz8Ep1jp5b602i5DqdkLBK9UcGXm3bpfSQdfn4/CXfQsB+RtgDEHIkZmADbpi9p
wMVL5sCZIRZH9sfm5eVS6h4WlXTHbCqdaBPIAufmN8yAnmDRpW+C+z0spUb61J9byy0n44/awVko
aBXI4CjK4l3VkZmIa1fZw4TphJgCjaCyuej2BRGlptdJlNtHjKGa2cFFNcWV7AYpuFp8wMlp7n8K
YMMnjo4gKvgw4MNlozyEUi4NocPYw18+n9OAw1JexD2Lni/dyuf3LnsGsERBVsJpIFLLg9oCn9Md
DxyLxPdhLsntH6SvNV1Hw/hzp06l1w1OXt+hch2/7mKIpUTSyhqTft2NS2+gunGoPaKPeSm7fSe6
A3DZxTZAD+r/VLzsx5wm6qv5ZQhxXCdSUVtT0cbNGMhAr2qpfGYWUR9/jbavhnJ5ULiPYNO8pxfF
MqM8/hPNRdrQwd2BvvmAItvoX9/fTx7Uc5S2XXVfx3r8v5M5Sc2CewM2mqs0NZKwIvmh78VPC1Dv
YcKHeFPhzmDsfjHnffQS7I8B/4bgE3eFkftHWEvdVbjoTgAJG17LSxsaaeA1Fd14mJtEvl/73g4O
jp7YDcsGMIu/4Sy0Wfx2Df+wSEHw5Oafuwl7O4QCIlUBYgQ3fOsaGddOoQn1iYuD/7AHpU8i4CYt
CzxCvx5X0bFP3dr/QvO390b+KWcxvIil4cCVDh5XFD+vvfa3lyvnFjKNlSZoliYtzx1vY/KH2I5B
z+XwC4aIwFDu8g/9g85pTHIEYpquiOnsVel5q4xHOJ780E42h3U7gqxCvKqC4kCKkfzRIMF+pOkC
+yGLg7Z9rNCQgXIBtbDI+6nHgiLj5BGEGPPNtRIFrokeQGAj1wNq9qKUI1KJsFa9syKHcvnoMjTa
jKiGN7R8wyLkuBjOie1QUbSevkra5q2/c+6wCAS89KMhqPKuXX2UGfa0vVYUnsyeBybvHTwFK7Tn
CUWkUGBq3mVsBeM+uIxr5QHSyrlJ31Yzgb227K9tAJUhT0imuz41Grj1qY335hVVpZFUJr3LDsPt
ykGsrfVhPkB1exCTvpQtkNMolt1T5rbWKEe2WbwIzP07N0bFitnokQh7kpR1a+ZzqaGEgS0ykKd4
nSaCPxWwSZHMx5ZlfSEnEzrfaioZDLReftmBnfTds8R7piZYGzsSNc9q4nJL3coOh2u/DeZOHp8w
dCcu0M70nS/Pj9Hz3QIa4iViQYDYkozYlInuhQ39Vhsw8glCCSMlhclM3uyEN2VtX399wxV/iFiF
JFln0erXnHKi9baW37wj5cbmND0yU1CVvyEn//lunoKc8p5j1p99C/qKai3i4OgycvNK9gY5kdo5
Iv6118vzdD+qv0tUmKYiD1u6bgoscdhRAAZpHZihTZvhWCx7bPKPo8bEwVbcM8v/ofQWTyRrUtI3
0BZeYfmZ0ortEunTiEbDTJAqvp8OR4wJTZ6nuDS4w8x/vvmsaRSvgA+WwPM6rhOufJSLO8h308wx
lBVseh35kwYwM/N7VTVeTzI9FvqJ9/Z96E42TtzzmZMatr8k4t/djgyCHNIp8LFjFB+oNtmcLUlM
w47zf/3Q3JlEGYwxVMl2M5rdehrx1MQc7iAKVp2wcgmpz7SxdoyEy4fI7e3hWvRBi37BTi5Z9LDD
kbvsmEZ7kfTw5F5dNn3FsX2HHSnlsJkfH19LGpoKKYAocMmbnvLdNMN4WjtdP9pzkt1X4/s/RSAr
isq9UTSEpeAQtOpH7yX+Pry8MrjhdH40AxuxQuVMZwUTXYhoCBL5X4gZJBFOmWaJ1gVlKyCkYpce
G91r0vF0l3xdbl3iMhxSqUQQ6C2kp+bit2JmMyFM/SvDeqU3JNgC03ac2EieAMHEdkSsTrcBqNya
UVxYT75vMwNmwYDVRIAbL+bYnUeIWsTTAXf2ymNuP62HA4nBtPo1HlQ4aAk7CSiVUPUrj4478oHB
T1DxnBBRV3RF2shTbhuTY5it7r5A8wcPWQ9208XNJbDLbTBdeTyytfoER2b+ROuSRwK9tPNQpLbn
TubEwH3NDDUhalJa+DIrlT3LWUbCFJ1srtS4j4onuc8rNNfkkOYAs/GXL1J1wp6yR5icXyeOSkhD
aAqdXq0meYnYXJaR0HAyIcZGXPblWOFv/zQD6cXMS2i2C+PxANjW+OfAqN8o1ubNqQZ69wX67S8h
RoJu6gpJXUG2XtDsao6e/DuUVFOGfRT+VhYIX4viUWUoVR6lVI0O++glj/M4KfifP2HkMINv6U2R
IP8PWK+zgMgLJWYepg1dBcmbJdaLzQ+MxVET49GyNLpL+RhstszIqvQcvmuk5kBaDsqdWgPtw4Er
SC5RVaI5xE0l8foIIRXnQnkQJANqqCt02O0kqUwBvYSzKPiukFq5bZRJP2B5/DYVId0Mrt5YvvI7
lY0LvOwAvQCwbPmwQayyxnWQY7hVHFTbv7lUtzB5WjEohtwQjPpgW5W6/9wW/ALxmwf6UqoHQI9B
07rw5HPqpR5mURIxLXuoxnInFUkgOcLiURc1LQZ3tFQRcIUSptTwdasVs+TrXhw6prVDmf/tAzcR
W3887DDHY6vXCZHjymeFSK1DGJbypgnVkbB4OeKP+Dqa5UcLgJ3YegmK14hYJv54SZmfw1JohUW/
cRdRZMY8stHiwDmixZe51+jJhkvjUBqy5yQc6F+2FQriVpbC2NyDQTh6yMwb+OwbZK3EwDdTx1l6
eMzzQgNkMHv76tOp7Mm37Ak9dafH/YtMsXGJtOmx3MmUxvHPSkaK+byO0zxAqNoObSptIHpOXZ4L
RTt5EqgsywxTWOuDsFGbG0ZulcmbnySvue9/PXg7WikOS4UI0ApBf//ttvDXMo52A+vJKYTKUnjD
I8B3vKRNHArthEpTjN2nZJSfPypGAm3g6aZ7ehE40YkTGFCi3EObJGWYT2wtJtzVMrPaCMTgCHLa
1RrvrYUcD0s6rzftmBHMjWWHRXHBL3hgcSfib5BA5YvT/mpvzp0MX1SGsjqHxOiTNQrOoKbivlsF
Vx9Rj5yy0gRoAUMWBV8bXJMz9S3UQv6vx6VK19AzPkz8T2Hq2SVhLnA+grvOk7RnABHkrWTwlfju
PbMuNab8Wgdk6+zRc2L2umciMRTP/oIlqhGDDkM3dW2eigNWJqsHwSbiQlSLNoMBMjzX0VllTXw5
QzsBzcJtTHePr3JOUTf/CctnQHGfYKAhiPpwqal19ginPuCmwIW5jhO42ARVZ39WLXTMkxDpf6Ol
d0IN2H6EtdjgBLsLzOVqpI9W6ZlaSD+hPfeAug5bG2H6dzOpNVczzfDQedD+I+FUT8CKEqVCpAe9
mGMwWMeX1cSk8FZ327rpi+ZFHAQDJX4PtKMCjlFtX9yp8ZqEbp7Zydun7ZhvCfawnYmzCKO4pCmm
5fxZk2tpKZP8Y/1o5s2f1+YAEWonDmXmnywQ/kske/f3jHyeXBviQSDvSyMepLdCpjLT/0b0ceYA
KuYNZo6aizIJrc4yEtYMlHRjKdyfGB9NTH1IEucNQlcpQI4nqf2h6Pa+g+lyJCOwsNxqA9eB1Cgx
t5GXrS2903fKBJgZEgY/CJEb5o6jxDd+IaxAohIOeeweRqJcv0/5Bqm4y1BLWo+cLVVs9/SSjwJV
FcYuayt0RPOpTWPlvxWJ4gRVggRR7rgdH+TI8tIZSZp8z9OaSD9HEBYS9Lj5nnZzU2MZwan/L9k9
9GsxZhNukSHpJmXEJLpKwnDXu0jCuLEBKAm0sfOTKb4CcwZUzbZugFifoKlAVnOAvC9UKD7JsWo/
UNcqA+7OhgqBTeMxhtqN/QBNLcwjTdwlV7emMglb2JxnN03swsKhkjwb72AGef9pVVuBr6321KEn
d8Ua0CHQnb+NkTT13q+dulQELLFbeo//MpD5RSs3sHl3GvwUXHtWJFtTnrSloORYVn4QWApE+5eX
I+/WbbQUyMWXFL2ufCr7Y3B7uAwpTtrDvUrf4Ms0LC7pyAJBqJ+qL+ehZWWliZZyfHXDVapOoo6L
NNFEMEDfg8SBq0VsJWXOxG/b7A7iBe/pmMykTUkF24ZapE8L2Upa3eiKxobXEKSVx8qZsJQtBU3r
bGoqnSlje+oEd3sAbkux7jpbzSJTpIDtFk//rWDFSatNjLGrmyRg8UL+M38/YydNbXWd7ZFfoXpn
f1CK2rDMTmZ6/IuZSB0ML+jWKFSZ3EDWnivY0TuXsDBaXUFaSViDLHC3AHktt9q7/3MoI1+1mrH6
onHiFov/iFt3+GM870EMDPKvhTNR3fQANIOYdIpv+svWoi5ZtcrMH7Ro8a0Ya4XYZUAP1Zh0kmV1
3CEg5Et0HkgbUVWRhknDgCD9IB/gDosqywt2SL4VH0Bj1ssFypuwMhjhCC6hF4NBvGvjn1sXzIO2
mfvPduhv9KnZhHgTFDHHStLuKH/LibVwbBU4A22hxxpxnD61Qhj0X5lBIr6wEJPF+sKXqfZYu0xa
xBh7VJN7q8OV46TSwAlkWkvQaXyZRr57GswKR+WzpbfVs94o76WlHzcdVfIixFfWRLVc+gCdkn9s
ZrYr/T5nggv9EmqnpLN2s7wOypxLYm8GpAVTakJ7gkG2gKPa+7oqgHdvpqqfh3flput9qzvQ8W9i
94Kz8Ei9J1uvx5BtKyHSqmDrDWtUFFl06il+vq1dDeYDJRE3p5ZgLAO+DWCKgfz6iuTNQV5Rg9Xd
An0sZOiGEBKIwk5NJbkRANp2YWpA7+s1pSyT8JD20isUVpnyq21U3RWNcCxcpygAsQ7YwJjxnJF9
EmAI/5PvHfXn7djv+FM4G8GnoQBcj2lksCxnzC9mXazTt6xkuqQpUw+xRYRBB8VIKZgG+fdWljjc
zMFAsWHsosA4Vrtcl40dul+SA6CGa4Rnlh+g/JPk65p91V+4O05CB0y4sdj6xSCU0VJlhZcSb6a8
/2kh3apdsii65rXAiz88QZ+by7A12yJXvCBIZcPxSWkrbXo2s3GlcQ4YFaofmu56TlFuuSGZEJ1V
D/K2mvJbzxQvl0ZI1Lp2FWvVZPIQF+21/berSMbSEgMV63OWoIGAPt0AUR3q6GTUN8vqaEihTvTT
BXj3WvL60PQjl1qBRXbctKGEJcOmxqQxBlVo6RmGx+lizwqCzKX5IGAExnbISEcndZ9Yv3p5H7g8
wSA8s57a9ILIqYM7la7EZsfT4DmyUbLoMb2IlmVgy/zJ+TU/WNL8hCQE7zR1pVUBEvA87cU75qBl
VYhiHT6KPVRnc+Smv0ILPCb+pBTZ5FsZ6syUnq9NTOU1trRcKEN4QWPMUBma0Sds1Z42/xqwi4DG
kOEyU/KiM/fY+d2cpI/aU96hxpvEoB2fpQzaV3QDR3jbHgtcpfnONktZeoZJZHHHJ8ETNRpll2GH
Y9QWqhqMn8fuUIQ5AgqePv9phhjvmaHRKEB11clU6uc/ul+/AyhPxuMOyk2ySwajOX8HK9yng69+
Hn6AdOwsZEuqguzWEErT9HHs73A/oIXUybIu4t3+FEL+3KbxukjIrCUq8snizWruIu3lbsg25L7F
CSRICsRCMH0K0g+hptQ00coJp+tpUPg/LMUGCQql6gBgS0gHDXr1N/ZXHXKrKev5YVn3M3+jVi6y
SQuBsVlgm7ee8KebkLMdSrt2X7Rbj/6O/bIbpcrbNMkpzSrAKaMarF7K7/gte3Z2Olpf/6PJnb5u
kpYRBY9sMu/FF2/dza895RoVgMqp82rMELgy9ufHpV6yUMx+j9hOrWFdV4G6To4Xgng+d6uOFcU5
6/usC79MGMSOzoAKmiG6eCJNYBwwwfOePMuv8nY+bpIqtfCZfTmgP9saru00PD5wfwCIn6wjLpWy
9YrGaF71HWg7CE1W4hvmQ0kIEWNzhcxSf31N1scNr8KJTJVSbbTFHoAxsESR4lMCLL8wcK3aFYWB
wRNuZW9xhy3xifQsE11pPtM1rlBpxYP+dPj0xIEr5uCyObupNsr6dWzTDhsvL51x1Ht8qWlaiIxO
Q0PXHOQ1d28wwRPj3qhfbCys5Z/MGdNanJrNIaqNReghS0qTYqavuUdSIXRl+BdqQimbyAnQ/7OX
X1s106s4gJ/iiXRMJ+qjIJxnkn9MzibgrWdNtK6STk5e+aAb52n4rbolCB8zlw39e2eR+GHYBuFr
8F8ubnougRJdSaFskJeMLeReEdh/hmwdvu2rlS4l8Yswfr7Wq6DKPv80mQ40k8RziJOJqN9uWKlX
tCGz2oDUj4jqIfeKFE8SFN3qDzZ/cb6HDZV5C7w8LmZXuwiCN02z3iOXeZvC9ZkPu10ogT7y2mEh
TVACuDeRK9vHv1UtHUev0i4D+NHlUvC4gPNNwxxpVA8i0X4bozJIC0RRrqlq3gyPZvqB4g59QfYW
4qRV+lPDMt3Fr/f2GE5oEb7T4JYACYdB7w92NMgNbF+Tig5lxiFqKaB3Sgp4Xu83cGCNcOMA3iNH
voxbS+dauFuKop4HzcCTtF9fDZ2FBkEOjfnScCMNfQJvoS20bbq5g0R37E+hBcShYT2FZ/Q+2Tkj
KPIE0Th4Wm3Y7enMppom8jfYdxA3jAOQh4Wox3NOZC1NOALgSL71URFU4Qi9nWYLBO7qN5aWM8Sa
eQYNZjJQoRqgHXfpaWkG+iwoOxP8wpl+eAPvuxKbJuzN0p2nuOeffZxAvTCDRg/dc3JBA6A+qoDs
jCH9SISks09MoihfOwBGe//Yt1fXJJLQxygwPXxIDF1w2IP8nza5MY+OxVpu7yzA8d5iA2PQlRLc
chJu6UWcmVCWWkmzbA4JtRlAZTL3khR0epxwF3Z7lY6yQB3tcsoGIiGimT/L0m7N2kAOqA6z5gix
/0ha/qsgZWZHT9WQVTlZGeL98SC+7uyvO5xjEsMCGdkwGXzpevfWl9bqku6y6dPK8sBgcGqTUnqZ
0wubbDOGv6O0EUOy2751Ny/5uhFFG7CZLWyWLUa2tZDIob6Vky+dKVoTJ2oTt4dvd3zSQNB9xZrA
DNBQ5K0uEUOTfYfq7LrgwC/DB3rOyntlVU25jOiENdgj0tmX8e5ZaRGiaLr89Pn47oSAUAQf1w06
TvrC7sh72CVog/aawuI0B+EtIv432lkrYbdii30N6yT7scWBiwSmSWrBrXpocEk+wlz4LtqoyTD3
I36ZkSnxvLAwnR4OAWfxMwFR2hbBWdX1HPn2SyUH0vzKuuR/wcT5y0FIFuWPcXM4ziu4kxomDhlX
6B3eSnltTv9QXSKBBkaCpSzryhNRKFmCrBmtk6PjiftrBTqAwcaHchHxeNr4zGKfxDtb+YlKvuK/
2XF4SNrZwU17UqHO2PvY4Rru+YA7NXcGk8EuIeb4+NDAz0bv15VH40vsaiLeJezsfTpZqCI/N+bt
TudnNPgfjGYjgL1NPlxi///8BI33/AUVWCBMVuMGXqWwKtb9r+LiJEWtWnTLgG8XQOvbL+rZNRww
jMf/X2/ij1Xk+EnmC9eAYl4X/YomARk9mqHf1oh5j8qB6duuFIbsdKQIUjq8t0sw2sHZHF5fca+s
BxLbi7RUpKvRshkZMWBlA0CIzJIPD+9DwgXkbQH4Nz92uRAc5UWpNs1iIHGqz4TUGLJSmw+0Vzm8
WTYsiywagKf6eSgAF3Bl+Ijt26v/Ez/JYBI5HEtlbfoKCX625gxj3/siRawuAt/euxC6ZYXVhYrO
fUXwAL3ksZgsavkV3jpSvG1Rlh38lEbsD6Op+tlbFcwU11vG5ItU3SO7r5ssUMYaWo/6HNHrUzME
A0TGTwk5Shen6VxOGAP+DbV2FQK+V9SdUmY8hT3PrAgpnXPQh7TroMBANmzWpvrCTtgWyducaZOf
Nr7bIDIbEQ+LPQFZSccz8ktpn02iJldkaDpQwfo2hGrfoJzEWVbuIHxwzbfLHWKlQ7aD4Y2ixYMj
vILoURv65t7J7bPK1v1U2GSvbXmGaX2VJLavObcQFQejNyONlUULCZaNH+CSIs9OfSp0NcM5UjMz
/OBjwN4b4rQIjOJa0djG+TWr7l0snX9ycqZdJY2nbjwV/q+0bvlEgPsVPnbblpb6AZp7zKS2NdEG
+Lk20wqE16qwyoFkvJ8+BbfSBRqH4zzA7UMd6z8jQ0YrkPLCtzA8CVnxzEBpyRPpZYw7Ess23d9C
V6u2o1vm93xk1IaPPMG7cppb8f2M4pQPMoNgDIGUsZCg/rMp/eCkgln/+wrmwypiUWD8n7pTqoj0
DGb/d4wy1ItPQ29e93wUzf7rpXdNmWrr99+pw+1ZcOPwpUuX7NN3u5DXvDMCx2nyyO40lhhrK+9I
MKq0Dv2HfEFLvO8lTX4eIbMbHkMbkr9DpNLL+OpCuywDik0TPVwzNVvTwV+9AXqYZUbFeYN2cWkN
z1RVbT2sHkW1Jv+LAEDgberRdElQD768pYpBtXrDBe50qx0hEH5liC07lEqqO9Nl0vzwzhgfcwGI
25UXZ8BKx3IbtKHZTr2/m3weEALvCTKkK0FU1Apk1dRbtwL8YVG3Ko5sg9U5BMVCKrVr83Oq0Qhz
WyZ5nTH5x5/jpbBQq3u4Qp3YOSTdSTLFB6qBFspfKr+mzkDjs3023TGObdoqVJSYJm/N+Ya9NLTk
+cb/m2MHhXpYIwEJea6pvzLFF1u8ziNtcbjEbW0ILX+g0RKZ6W3faq61ShsLkS2aUm3upv+mDr9l
YLIuFwGpRBW0N2l5UskwPoW5fSmzN07YRf+GW+c5hfhblPJfJslQUBGrLv/E/buSR1HzGAGwhP9X
bONkbtflNbEhGxX1ebjJ4CcWETqolbnsC7vEozWGM9zlDzNYHSsmWqDKlxwXcz3QyWE3env4lIDO
THiD7SnopsslNOwOlzDhD45xCAXpVCyrZvh5hRek147eqXpA6rN785BJbex4T9UGRfZr5kccsBqP
CcjcHkThTQJDXfumSe39m4nwAtANlPIyXBxyvhYTJr2sZP/qt04GO7L9ZeLwAOGJZ35jFXTEmqLQ
VlgX0+WIoyQJ2ohFYLx5M00OTuoQBbs1gU5kce3XRBw6fKpmLwVUqMz67A3v5+SdRjvWC9BQyTkN
WcIqMtLKs6/+Mzhm09Roqfvz2bBLHpyXqqvMGWppaB3IqrxVTMj9W9X6NdFkXRdkrBxp/AJu2eJO
0p5U+bBCxrHIPuzG8SDTO+Q92v6+XhAGoUAroPxnvZY7GPZEZFhLn8bNqtP/l7jviuu+o+wqNHdu
FhX5m+4HigVsfAxBUEWZMpG7mOifcNLvbjriSa7Ki9FAv/PC6b9LM5Bs+FE7oGK2yJJL/12Y5Oer
SnX3XcZuFON4TyHaaTRYWgmoo7pX5+WsohA0fFcPcHI+SabpjIlM1vqrPqiN7FazngeLLgQDiRf2
2MDSMecyhXP2tSG52q+bZavRFeIbsbnf+nIwdUDFMpWv47O7kEhZyJZKgBUThNCY2+WNG5Qa0MQR
a2Z8IejkK5xVauNp3VL0Pfb/uIqTAmLgAGfGiRM/5QqMzTwbK8fjatRY2eVncedQnukpQ0x/Xxhw
n6uhc/J1JxCpjYMOZ09g6Da6AN5vkViujewVnseuuvsgpg6wJuP1JatlsgxlE+DZWn8mNU7RdDbK
TG4oQGBD7j5GsO/O03qAmxZQ7pZ22XX5rNT6bVCLM1d21W0seC2QQui9o+EnR9ImDkrBUD6byi0a
DOGqqZtukbmqkfD20SJU3n5+A2GBudjE0DqT9T8ZI1fql+spYCFqb4mvhIG/K0KKexd+67DaZVnJ
vIAM+xA6OonwCn00o9FQJXLb8Q5QYeRQ/LffrctY1FQSq1df/b78vNBckp8fcaoZjqBdUMKpka1Q
l58s8m2/xk/AWsKM13u139rtFUcTdLZ6FYalgCdKzmkN+chAvgkPeFj3l7NHYiaUk/WqLrN7QPkJ
QaBtePK/tLHOoV2wAkpMqPbVK1He8wzOK1GbETa1qtaBTXCWsVEs5Zxl66SBFCc3qe+S+mwZ/tlM
FMAhfXIkNKBuALtXB1fb0ag/lgbq0gJRPmsXGQWR7cFkQJ4m6+lxgHDC0DLeCQQLhoXfShlxmjWs
MOOWWRS/pMZMY50rCX6gRXrYKcOM7iqbMRqq664hbGaSsM0ZRDEN5rs0pSCjP+nhIV7OylMRn9ys
rsMH0ARp4L2pgmaZQESSJyDkhND9vuOY+cM/FyCVGsPa9HnIP5QtHw3zL4fckWff3sLHq7CbaYf2
WXLsQuB6un8NiPRfEqr2pVMac9faRW2k66f96joJ6n10SYowU01Ea8sjFPADps/oTTBS4N/GPgp/
YW7ntxQLffa5npYsmVOUr3/eVxVR6JsqMQap/a8f4wJjWojZ13J1LFKJyE13T6IeYJPkrUUt3ZXZ
tYD3qn02WX/3Bad233tkM/3SB2yquiaGmJy6g/3v+w2/xZgEOZFse1ctiB/7GKxQaLnuwRmOXfCT
A72iezcRI/eICtmKPwKZ9XA+XCj75LWRdg2cKLOGU2NlCoz7mPzqlMmL5mqK2peK+STGGmcs2iKF
U9CDDGeUUkggGyvH17SAurowFwxsusBQ5fLGRaLUVfDEeyodYLTf689I2+vz7OuqRj8PRBpiM5ug
Nxai8xRayFuWw47XvypBIWM3CDyk3D6NXN62xPpUmU9HZqg4cvSWb1U3UN7avTblpI+M+78+B7vb
MhHEG5FgYFc/egnKRJr3kZbqw/PYcCe6vF68TgPO9SyF0qRL9o/HZjKBZkWYSaWSoy8wRahoou9T
atH292qhKIGaBGClswwM0Yc9CDEJklW6SKp0Rpg6e5TPYQ2qHIvZpJFLxUEcN/N0z92GWtKm/dYh
NLjv+68epFl8GK1Jel6wPkp4DjtJNF+cUnPJr+1Rba3HsXXh9tpd9gRdrYuQq/yf8MRlM6atyfwQ
zcMbhIc00mffcNLc1z+M+FPCAziYVLHpqz0dQpa3MNWsbvpWEkdEw4lcqXSOpaQhfKL1aNn+s+GL
IKdQwOxXVy8EqBT7qgvhMn9xwOXvh8lMVB/cZGrlokPLxQfKTS+GGIP1y2pNV0teUyVhW3dB25Mx
6tvjGenYLY9IZzUBNJ/uLkJHWOoP6XVj7EZEOXqapxvWtYEdP3gWZy1gjdnnmdlHss310KMATK3k
Q3g3v+UrUTV5kvdaBtjWlA/ThdHvA8HxYwt1S8jEU4+wnpywTTYUFLFs52xTaCUKu5+dLTnsIkdv
ZJPHBzOrF+Vyt3gsHZthQ8a3G3weAvc/khkUo6RJQoeTwZIbsIf5KkJB3gAUeMOt6aVfc7a2bCnY
AehhLZMXSgHoYyKBr4/stA/in5fXwg7Wr8fZ7+8hU8GvAQg9osGo/z0RPcI1C5dKITtSkUnEazJS
yoiXgDqmaPBJX/nQyCITu9WFZjYvL4EP4K4BN/jh1LrWNri9Mzryc9WMxYF0VVy22q899H/3dkJ6
IPSs+62P3TMGCyCkosusO+/w87YH3lGhQKWAWaUTTiilpEL4UxTB5+t2nExTK5gLGfaBS6rQKzDk
J3KAs2tF7fnC0ptiicibmSFmKLfdNhq/DHDeSTvr9ORgn/7ZKkKKXyuq/BNcp/LQ67eiGymCwAgf
p4FSsddt6dVGy0tW4dbqw8Qc8l3iu3rhVGc/R7CYFgw9CbUP64y93LgjtWfGLDTDbNNKvo9YrlSu
kQiqS0aIBAxqMg6rkNseC0XeTDvCuoVrDVgCYboEGV1XN8TnoXICG8y0fV6hmpuErzomKtP8SJa7
net/m5hcz95A55nAXSsCQrFItBH8GOy8jJYzlG3Nt5XNv6FtgcmAgJU5T2LjvP7lRNIVFyKYAY46
q9hRCRR18vo1axuS6+vleY3mx7YKc+m/R+YbmlqRi48Y0uOFIqW/KgO4qFIOw7k8vsoEkG47qX8Q
44L5m4KDyLI66RBlyPoYiD4VcwZqIoJvykSVOroJRTEgtEv4b7YU4RIrbjOg2xWi/i6Az8ZJQHZ+
CpYxJhhu+pEwIgG1QszxMcItycLhjjV2VckjcyWNYnr55JS1U4F0JidvTLt6ydBKQKLgbR+ZnZvT
J9Rld2WQPx47RnHsC5lvYESa1NxP1PKbP4FsI+8MQ3sUA4S/hW8C0fA5zE0nCtYWasj2WyATu2oc
IHPHx4kb1f3KP/qd9VDADZdCknZzsbXztJ0vYmclgiKwgD8QXHgvI9YL5MRBQ316XI+B4JGLDSxI
L7c5eHGMFv2pr4myATZp1cGt/wdI3xlVfJ/EP983V4C0czuHvmgMttIc0xeGNvpenxy07KFr9Ad/
MJuON9nErXW/sTjABOVtz0pDNnto00uUZf7xn/iVecbO9Ry4hv67ie2VepWVb+9L8SMkKiUKJQAZ
pSRBAeE9tsRHJKqioLn6170TOW2wtk3h7xn6LBtPxVrsQ2ZlQME+FRqaDxVN3wkv8OVNRcxlimt1
wVarthByUG9oI0bVo42U43KVrH9/bnupBGrLAJVru+zyZCSmcCvbC9Z4+KXsPTEe7vx0yCgJ1OrI
XpLFv5kDRiFxnf7UbzHZo9bOAnbSqahl5wotELHS/wF3L7+HSq8Bfgc5KJ9uaZa/16QCJqrp8MwJ
YXYI9fH1t69cXj4u+4mIepnNkaDDX18tYZ8NecEiVOf8mE2FTYUejJkFfd+NOJChCKuR7FGM1QtL
fttlZo4GGYaZmw2XEBn2JUlDXOLxlvVrMWbFeKS/YNd4PQrPy3THVlMbP/mhm/pVUFB7/ui01Hu/
7Hy8lVQpBhp+MQq6UGdEVok2MTI8iA7wMGmcU/UIRnYUdPNB3oo2oUfEKiXhIaLr+NIJ5oKABKBr
vEUOclyaFvaAW26MUf6LKYgpwNA0V0hLDCKDDp8Ly0TrF6p+B979RIOlLI6jsJIgOMLOuP3V/mdS
uHR+8iwrqBxXLSrxymzaPUsMDQfXPVXAb2DpDW7hl/4tZCq4B1KvDQcozNtNShPBLcp2+TcAqveg
DdrtiIMJbBSGuFZZnAn7z99esPbBd04CBIpiW3RixwHXrNelVNaWM8B6dEM7ICgybKbywigBFmJv
Y4iXUP1knrwwF6ZUM6GYAOCIriLCZ/aMOYW9D2Z7xun92gdpAn437TH1FbLx6TpxgdEnLbE4/+Qy
lVAUuMXTfckFrlIOvdqkIM0JzpEt+CvD2t5Lpy7Fzfgso3InnRcIJgAUHTTUcDf6kq08Y1rqsGNZ
KEk9We5M5Eg5LOO3jTA1rdGmG4pxLNZufNdailgsQyWwx4zB9vW0wnztxdnPreFLMOlHxt8Hcc4+
lvjctU0p5LhAEQiUejyEABShYGQsqi8Kn8SDxoxf4X0YULWU+u5hD/iNYO2aXECcnGg7cIDT3NEC
ZAy3hGA7N9rFItsnSgEyxoCiep2pUrsavOR9RYgVYxfuHyqvLRZDFajf1S4re36njxWySrKLM91W
urLlOH6W/exb3LDcOZhh4G8y4MMblswcIakokZzGraT3jb63efdSinhEplD0CsfiUDBxde+fKL71
AepqxgkZb4GmVwqfUYkuNndjbL4Lj4jPt51z4ZnRAujWaxe2haTkuiTtA4mWmfX6n39eORa9pvZW
lJI/vXumjrYWqZMCi+1gkaGtAA+38VLXGzBAbLgHTm6xBHe0eSJl+3/9olK4awpcCwDYqlKmp/vL
BzUW6mCvIbewVQZMMKUctVdCoo4yW7hNr+a4WmbqI9vYk8uKTD63h4rhoZYRf2Yl7A8YnGIudcl/
sxAKJwljwh089/ewPV2ffUsKurHK7iX/vRfSRklotySaMNktOekswpHfgNeSmJKrVI1HsLmvu1Dm
VPYetvS8+xrBd5cyUOJueEXM++PA6bTNalanQyOUq5aK47dnn/0r+bR9JEUazjQm9AvFaPP+ARpH
uGPDR+ssZwRhYhK5tKyfqwpCq22B/VXGjU8XSSxmwg17qETKlZFHpzRkzH5HyDiR9OJTYe5qVvMP
ivOUWlticNsrZoX+GU1PSIB2ArZT3iwPw4rnPvGG2bAUXXinIX9/q+zePUyFpkp1IbeDVSZbT1o0
4mWe9n1ayC2dquW8fODqWiQoSl2O+7YcJ3pNIc0VpfoR6gaQpoyxshsnOMMPYGn4tEeJ25KAVMzK
n7Az+sBMA6ZhS7pW4bN3iW8F/hBczREj/++njtDS0qguMUq97UWxvfXfJ+uXOmdr8lskLR+jrYnW
nVuAV2B6Z4f4vDB63P8UO/llwDOsCzbAqBjclFNabI+VWWCe1pdKnk4cy7cqhrQFZcicToIATXvD
cqm7jy0dfHFdwYCfIjDRVRCEeTZ+ap6f/6JeA1kJ9ZXuxy/F0rHYFtf0CRTFPKuaZbaJUffGlaLX
7tOnq7vCHU6j2OpfsjmsvwE2G8pycuLX2ul5TzejXhA5eDOtckHkZIf/Pbru0wNFQKXRQsFAAdih
jbEmpUtF0/DOuNZ6JiBwZgGs5EcD4i+2IChOUOIQGXg+hfLY6Vuh8hQNUE2JzbegPMugUZ8hGCcX
pmCZb6xWwqwnvZAHud7kBgcry9Z80jixtUutrsYNy1Sb+RksFCHuD2appyfICSC8vuLoAxsXGgaI
v6uTiVlWItZPv1KSeir2x0ji0sHksMdlmXgcZvNbGLIBZf3EQ4Wdj6Q6ZweBotkfShQFxPpl6gan
+AVWX5J+j7/LEPv7pKGGh610fuQaoA4cYF/x9QJEXmq4r04zbaVWlqtbYCdVpx3clMDDuWwKnYGH
qqOuhUYUkEJd/Mdvp/RZsryRGboBX5yqyfUwRDNEUGxGBAiZygG2tqJC72jTTmVlx1g4f9h18qzW
64Bz4gdmBRip63BOqxsSXXkJI5qfa36JXrzSscDYDnsFH2CMSe/Cl5l/1uNKqahwTxO51DwxCmZa
nOQZgGpbfD0TdWiQliwUUIyfTOJSvuYITzhlzilaRrM5g63yBpVlgFiMy9byqOXDMS7tyI8phap1
sxx1Z3ZfEbyWzKBmXSnN73uHhLSpod0arnpMKs6Wn0Wy95lciiBzeUFZvElUU3wnhFyDdZaoKksR
4xmJ6NJaDj5gR4Jhydtfo5cORZ4glhNocr207ubDz57+gd/fN2HNAaBnONkJ1YzP4lU7qd95HTu8
dgirRdotBWFSmwBrk+nlfLRPV13z8V/4dYuLLQxvwqPA2cGs36Fsyx9s34lNght7D1SUhhyTSqMe
CqEt3GLJezoEutpoqlmKvr9GshhpK95AjAy6JfDccLt6njjfelLx6Gd5K8oV6ehGg3L1/0u5cMPY
uuKNBW232n9pMBFrVBb4Gmu+fOJVXn/3G5qGFxsuzfbIyd+FYgraxdKR0McU9l5t6yM+Sg0IGySh
KGX5AQ8Yv8FJjVx6KPMSqphvnR0mu3GYoZI5whVUvNHq9NBm/gxUA1yKgChEQaoBipK//qYDp6x6
xezSbIUgQZpRGx0dnL7VFOo6u/lvIvgpZfSVJwrvVqP6S5gq1fLNZi8sdE3vPH2pBItzf4WlHxwL
0DnapEkAIbI4OUZb/zKydUHS0yXREbokADWSepxYSOHoT7+c52PTHPaEGk5B+3gGusTXIuyDKk+r
wQ1Mfu2rqYDisMxL9yIfIlSJBK+8UQW0GQNi6aH7fUI7+JqmJ/ni1JsTiwo8CQYogLnABdrULRZ1
lDdkSqYu/oW75RNuxqZ3O85PKK3VJGrnSiqKeHvNqyHJ2yCrhyGWpIqItrYU+4tdSpC3sNDBTmxk
euAKqf15E/LWr2Ih9LmItxUMyZ1hkAlNKBUWw1z6D9bCJLUzdGrpWkch7DY1PnYgtq0qRS6pbPoS
Mqy5SLyshjYyBISBz9Bg9xAKaOr4Sqqfjj0tjItWjxIDTbCaXOfj6xUzrryUKKQ9FCgKK2ND63MP
qbrAiPdTabI2fQJR/gwNFno1VjnCpdl4ITmANtJvDqF0o0e5ULnN4JMytpLzvu1ia6pqaRPXCotK
8NRi3GsxFEkuSHzFRHGAd5GdxWlOZovOlJUmyOVNA+sQDjSw2cbIaiUx1W+HjcoaM2ozPGpgBuii
pEwjybXyrmq+PTt9MQo00mXINbGGeyBqzF1Nx8I53Y/yms98P6aKy9r6pX+9CsSchC9+s46kKhco
co57/GL2K98OoO/7vvC6Mq0rexyBFsXYYBZrQeRaph8oJDOmlKMMTufKBYvD9p7cHbcDqUVSGWm2
hIVjr94LyzfOZoJljQ1ay4OwMu0EMF+EbobeAO8LQxrxWKc5mGVe9nfirNBH3EnqN76grZHCUu8e
pXFaDXndThJxqCLdT+LHLrP79iYwvO3HfoumeBXgDWl5LaZkj43xqdxIyElM0NMgBfh5zwtsYMRD
S24vLRvBOr+OemX+zcXLSTtBtfMTO+vnZBzU3GBNUnnAX7T+mnRzTsDy0aGEdKQLMO7ABo/cxSOY
TrtCOA4y9t/Y2nJFCj5R+SDsjDRJF/q0XiXfxsZKu4DyjEW0V6LAK4X2LT1sEUjwY4GGOReB38xx
Zz6ILwUnJHwEOd5IT9wBMawZbZXh6g/h3BG3PXqMKAyQTuL4QE+94pgBYN52G7JJp7CWtnz2+c59
q55oVIpRRBRp2/jv7ERJF34uNOiEmOPsEOlb5W72xbYDeLP16MtVQTDsN1ZWlt62uraHnV/d4vge
EcX7TFkiZE6XqD/YSyxjcvQOEWfhhx8r1X1vwK9gB0wr4SOuAokVVI0ega+iAD41o7COarURisu6
3BRxmVDCVWtr6z7vp+OinM8fXSJkq3x+XjafxI/uEt/qDJu+0+2EVV+0vGZNL54KrDY19FJotbpT
tHGZuimUVrvcZBA3laQQuCf8P9JBKniPRag0p8J6tMowPwjKgEP5ikI4tBaDmJD/pjlsNvR+um/k
5UfyciMhx9mq7q5ix0I4Q6/+qvnigwTQcXSe5VH5oEwiJLl3uc7ThJcTFg3OJkbPCGxRdOJ2yxDk
+X/O+ZP+ip5wLJc0pDfkLhegmKS5Gr1XOAcN527cl3wMVgGNV34Fg42yu43JYv85eW4/aQ4gurv3
U468VMIQnYkR/OA8wuHX8oyXAqCLblHvVJqZWxSg2mgiw/2rq+9ecSFT3rgI8bykhutrozmQbSTG
8De5Gvnny+qAmuOGRKlPIuWAsZHk1RlLXGAaYgE25DNjMKgXzgh/mS7VFN3ObPxY/vjcw4TXiouT
cEbwuNEIO33SJRXrqRsJJuVM4hxLhosT4EUY6SAvkJr+N44KGlModYRdYuvNLbfgJlSgVstAqb39
wp+trEHo6ztDH97nmtbD1azK730zmLEnwNtucojpINU3OMYOt9GvsOxKcPN2d59b4Q3qQUqSf8Fr
8dfa1LVGpgd2HScldxNJcWLTYNCUsZorgI0CW8eMfFN6YgPLC8v2u3P5gKMO6sPybha8IpvjCzO2
WygtSyBYvvsT9SeXClObUitlBINTHmLd5UFtW8g7Qqc95e9F4PIIwPECtkk5ezVpOCKirFFmH44i
9n5NjuJZsNmAx/AxLq9/pKEKCKPhl3Wr+AmLJwwubhANvineKqerg/AZeULhupOP8RlB26IzwFqd
qBBKxoL9/bEvpAecJugocrKCPPm1T3vDpag2oY+lR0s0sXCo+sy52Wu8X64iLpyf6Ni5KT23L23B
y0TBZBDKHsbwi4WZ3GbI/Ik5I3pDx1bwoQ5Jx5Rj5UVQ8zhKLlGTRTBnahsy3ElbIkAQRq1Y+RuM
a7FWx4Si7sUsB3gJavr5ADz5TP76zYHNJQyfXAkGq5XFpsznxPI6w1NziSsuFt7T+a4jUJGuDtqE
8YdMtOpPFZE6raCov862O+EcH+98mLaggSzDFG/5i3RmZ0EauLLlN7GYFBYIfEcu7gPeVFAI50nD
8H40RmTRtGu8VYwOD15sWO7gLqXni1ieQxh346WQS4Rg6kzhE1hwCUsxGC/3z32+gu1ZsG15vVO2
5mb17U5lciT/PgmsFMbSbecxUdBGKro+saq8pC3MWr+xH24zup+T8dVHhUuquLhxQwQk7pEY9JH3
y6GdEb/jYzIutKnXndAhFBg5QJXPKmsxck2ps3R2C3o3mhGzcFpYXh7aZR32QSDkoNlojxPoyy48
8kXFdmsPuQ+k//siqRnNZnK3mASO7AOig3yD9lL30k5nfJIZfzbUFOY6UVr3VnrL51J0M19OlkpV
T6zRtBwZkUIYTaFxBTWZfwMyMW45pOFaYKKPoorFWVXGETmqqr0qv5C/i6I5QZztrChFZy7nh1ip
o+CXr5p0eFTe3WD2P+lvj29igxBs5plIrEQ4yo+ba1hzsRCsXw6VP7VNyMUA0oAcmBvQY0X8zZn7
z9DOxejVO5QAViuUFEEX1yGEorjJSb8DHr/VtzMKHHR1WGFhwi3Vf4kPekcYB2tRmbc5gKHhiOMp
St+UHgIN72sSV9EQccIXQAiHCGaiBKgk4qNa0IbdZrJHUdZv9BLia8WhP865u9t+szq+/F8CMw9+
VUuHCC5BfGo6R3qnNkSL9fYqmFBS+ph2W9dtYU7vwMjoGK+C4C6PLWsK4A+qWL8fp0Bys4S5P8wc
rRk3ZGDsMAmKQL5dA2WpBU7n3bRNCQg3o4TVafMD0WIhX93W5ikCYaZ+UuPbqjHoMX93q1X4Abjc
RKF5LakaRdsmzbjDo4A/b/jt2S4M+N1zx3BR8B0ihWB1363/ThvHYWz1k2kunJ6JmJObWc67sxkW
Eb8OiIBZKZK5rgeQE0i5uSRi7WQTUzFKXO3igzXyn26eRgdlfql2ZJ/e/VZtSPG/VWBuJ7UYw1KS
tRzbUKzpii5tjoXZrDmG8nAfD9W3l7Enq5jQH5QIcT5OOmMlaTtsXCOHoADsI5iLM+wnVcUuXJAc
oAGGtHaV2hhp/AqFQ6hVamfBmpSYOuTQ6kwKwKpEhLOn9hW2ngb62s2cbfn9gWj6urOPJ6+s3wPP
R/cCFcv8nKR1SJSQFxJ2FdXsXUTMeMMsnnPahXF+H0K2diL+U7nHApnuRJc1FrzdnW8j9A1ubTuN
PIvaBj79Lg5O92wCgBje8h/txY8OKARzvNZMwQHwrgNwPQ/XXB9dK9JBZL08UVJ+OlQUFR4iyegx
0pZcxCX45wc5YkNQJXlMheeDfKc28xWyufPdTRgA3DAfbMHfbT4QK2lJpJjJ7osscCwx145dtXUK
zTbbUL+tupYkruBP3+Lkn42KEBHshxKSfcuAZhu1uygcdnGy7wNb+8p6CPMzr9J0Tif/NVeMpe50
5dB5GXdfekGxyJKMTNKe1RhjkfFvQ34b5ubdVcpO5fAzbkQnTV4f9G5bE0tXI0c/oiEUItLRJZiw
sIZJ6oPleLJdn/41cJxhhuaOBdqeaLVyNrd9Njrdzf0nyZaKfZf5CEAMJNU+HxrLue2BcOWDKf+E
hI+UhV0Z3AT6SglgLtOPpVa/AuReQLFPuU5F/gcLu9fpmW0UXW5b/E1mYSKe+8nzZxPYIsyoQDDz
9ew/vYwIWA7c1E3kyg51LmlblXvyc6g3OnzKJ/PJb6r2cU3SbzBPNYE2wQHEAAMzr57AVAOtpqem
t9r8EO0bVmXhPcDLNEoOT6/VGkhEHbs7++FUvDz0DYlNrZbXAZ8uhVGtckpgYTpRnbRQ9qzSYonr
Oxbm5qLhUbfDFR2+tplqT+bf24LVnxmHj09zByo2d2dvqnJui3GnYPnJGYu2YUANqzFANvPFz400
QJdmRuwubv7XFmfGeX9Wq8gMPCfoL4J0eLEo6Ay7oj5nyIk7jWSMWI2vceh/Rl0PTbitUgyUnzV1
i9iW1ToZWvxP5vNFwXMn1Zr9SqqyN7yDKWUEeTr713fCo9y2nNtqApfBwDF9JqLHuvANx7MbWCsG
eF0dRahnqnpLQrS807ofryYt17VH2AdLqnGxnCit+U2TCtpniuOkLFXE/oh1EpH2ndNf/h6/VwEq
rFhdLZk5WHzp6MfisSn0WTD9DZbAHQ2weYC8PYNnGCY3X6//3NoZe3je4CJ2bqdxM8bNIEAXNLd6
NpZ4cdd/SjVnimmjdcMc1+QFAndot6rTPQHdSnTE7BHkk73LBAWd4hm4Lbdx290iH7anisPVh1RK
fcKV1FOzfXeuQRhJP2EJ2NMYGF7TPI7JHh39B3jzZTtXYHQn76LWGVZeDSocDX3sjxU0+uKVz7Mu
us9Nz5GxhnRmzCtn9J/QT57txa8HFFFVaIqbRjTIGhk6bh3pfUP9pS+ci/hvQFb6ujuy6WqIpfp/
n8R2usYMq3TCE+vkXSujonb5QPSBTQgqQwFJ4T+/39+Igj4hJhMzTc8Om3QNII0aequxd40CQcu7
Qf5/s7xNGveJzQipDpWfICnYN2Pd3v33lDzYTn8g/9Jx92lFzYMV7TriNsVd0VeCJFCSjx3G4uRQ
2MsZL8Z9hUabqUjXge4BXP4+NltxDUNbKHH2dUjKitdeqOg3ft3YPSZ8dWWiYMtDl00KFr+H0SlX
ZNY2A+n101D3xJITDfzzbF/V9bdYiTFDIvhiFYtzCiQGoED+t8jjjT4us3Q+Ugp91wCfmwXaR+Yv
N/9QQ4i4WtfODSzxFQybiUnn8rFewFukmCoa9/ErRgBImEkTLxDhgZ20jpIf9NvkS1etE1x5z5cT
xZfCYfAww+XNQhHvWn/h2EXupm6Xxgc244ON7u8SYL4JRixM0qXu+IO9tcouFNCEAb0uc8VI+oCe
/cNJVZY9E7rqzE5lI32w2NLFOsmT4OczTynyKzD4fvtMnR+dyv9MvEsM8Y900gOS7mqhEs6aaMBy
9YOrkqA6Oc0knnP+olz+9ebUvxmQmi8Xl7b8/0Uuh3b1mV1ASuT+W8dNR1B26EF6a+lHFoQ6yCPq
Rr7jTNZoObGzk6wobkm8sskoaZe9G615hBkWgErUYHvNTSkffqINa/JczQ3GlkkNNgUEMMw0fHMa
aCWVze6KQ61DWfc1iMtpPlmZdkAopnNc5gvsDgvwRvUeL0GsWFaVkksEql6g3GhW1E8+zGXpBViv
kVKJYx3tFM4XaZQ6W0BK4UzfzhaPDGj4jDhBOHG8wWsHx055cvCfpWE5M7H3/CeRIBcjkKtHWw9m
G3LZeAvE2HbXnpfxjF5kP3UQTxCvGLcD0Fa+2vCWghyOwEM+JGOkkyu5PYT9UHpKzUaJesjZEVbq
7cOdAMszEu3GUBUpunahpOn4IyYtFbRD4Ionf4qHj4gGxBPMgfailkXPG7kN8LFZl14KeCyy4Byh
dSuYF/Egao/0arviLvrlvUr3wqZcfeW1Bm/VVdLvKHz2KwmkZRMsKQ558yGtQvcldBDxqk02gUug
o4mgBYhVEc37Y82peAwiSQ7iKn/9GIoKRkWCQyfXUptTxkoMVjTdjSLwHKce91um2cTPB/YN5ysa
xBtAxfGriQldsTpQ9MZTOif2ZMQYprNlFmVwIK1zTdQuYbQB/mF/VRS700oJjgZeX7JO2iOJHqMY
MErJuszy6bvXjVHSo7jaarnSy90pNk9EJjHtUqVc1LG+2OXRoPy1+PLMik/Ha210SlrFz3C9TI/X
8NN4r6jlP7MLvlBNTUVwRfDiqNtBYobf09PPUOAs89J+0oRSqRhcBou4bFgVyVaKwwQ6FLTU6KB+
CRLDmhSk1zL8S4nZpHl4p1ZQKJDH5e49iliPigGm+Yzo2E50uHjaI9QqpMoKJP3xmtpHWQUVAkQv
cM87YFIK0TRe66p0UZJSeVA5lXzPASakJq9BYryxikjQygV+8ywMa9Bmch3bjI8HMhmrQzjzeTAp
q/En1yNKNQjZg92V2uncl0J31N/Hk2m+Ht3BNHD4Gg1MZycpTiFVNR46x5WY5WllabwPVhgARdVQ
ec1jMeBFok5YfLmmIcluIUMEJJ7JcuiZx07Oyrm2/baQ1rArNuB/Z2MOxobFlK7pHqYvAmygZtP0
PY0x+/qlHzpcC6tEOGXd4rzMtYuhAkS4Zh+AbGARdV6WyHiJMEzE75CCI0yi+ZcjXeJZX8uEo/AR
kVQY8FQhrRiIzStvFm198JC7HSqyFVRlWUljhJGAizw9bCX9y41/eouwYJV028Lbrg02BE69IhgF
TjgncpmBQ74aF/yo3ufSeJStnX8Er+a0LyhDbJ+h5W54JfTRozCJNZ/8sAX3AKe45nlgfOxo+exW
r9hwD/NPSdJXQ+Rg83grg/nZgr7B75mNvcIUVMZ01+hLfEktrKxkOuLX5UwIx7vqt9xXp9KqZjz6
2x93SslZk4rV8/iG1JA3u3wqa5UfGkuna6qBeRHu7/+eLNDsUy3gOWBzboOsGiVTYFBp/hR8lkZ2
hHaQtSd8HwOVP8VAybCNZ4Lxhzx49Z+i9QzYML3SfSwPYeIhDVnYrJ83EMtFigs9mJqAM7pYA/al
HYIeTZwXNHkMnji3saaqN9i1Lt43RYRVcQivNZwzEdbcNSTxmkBj1LGX8Ti+V0qK0N+k5K6imstD
9EfjBccdkxwgJFb/PA0VKItCKdDi0SM5VAXTaDPtDK4qYA8ld3gooT7MY9ZrZH5aSGU+kM6PAlnn
WlFUyq5quWqR0XuoOQzHQqi9AQiFx+Vb4jkeial3H+vFH1wBi2M6yYy8nBrA8RvPgokImcmGXozT
ttzsIyXvIzvPTzdrsExa0uZ6P79+YN31o1L6ch15zLoOMo1EAfQk1CNHZ1kYXqgO2rvo4TQmVBwN
tHDcTdkStre3+32twOAIcc2arh6t8L5P1Ye9O0ibwrjFp13ZsBu71qGTNbiogNdnZ0WZDs9dxocp
RZY7gfeRvkaMPfGOCPSzFPTiiB27fz1ilab5Zh8Yc87NtOJNYEmN9ZySxxjauuOL4rPnIMRXfRuF
nhzZJwq/iWlixBz3D4yJOc5xIHsuUBadJUmYqWkDJeMPoeRBQtk4EZ8UfB/F9imUjnjsc7TEOeES
lH+tOaEIMa4dcrM0MJeONbmOgDIYBSIEZ8q48pZHWHZ5801soaUVwSmxdszqlya2ZMuhTFobTDHF
L6pbIwKeKZ6qn9IGDmDqT5eOgxyypNcaw17UmlkhSK3251JT5Rq57GB+XpUJE60ayJTdTilCZpgO
cv2MWktRDpWRfawcqEu/OuOEkJBTyj8sMKuI7Yg+MsswJLheosYBGCF/adpQKG8tnqBpWpsYuqR+
IHicRM+jLBnVA0N6UsIidJiz68joCfNX+IiPUKzFF9kE0prRaYch3uLqLsc7BRmKdzc/trLoBXEq
hZXoTU049XoCzCgwGWCCvaxjMY3oXdyt5XoDKJBR6rD22kBrJtTygPnePny8WbkL4QsVSPet8NXR
1n6Mls7ejmCJUkNdA38UXhIM8hd4NqcbokTSecJEIoLx503tGlottZb8mrQtQyMJT8zI4z9gwIr/
m5NgE70QULBnE2yEHBoRYxNzmq1nO8+NZwpT6yDB16jPC/+5A/wxYWQCO0GZttDrbDtqY3mC6gTI
bGVpu1UCi83f0rde1gG16O/EvjYMOdaC72NOKNPaHp5PTA7d5/sk3CQliAOhqM/li1gFiZ55yqCE
7nsQmr3tpGfgpHUe8+HcHc6rw+7yAsSKeSfkcu6TVZy9+lrQnLlgg1D02lkmD1fl12Gy0ls59MO0
qZ7q40pYQaT2i+7Rsam7L24TE3Hksl+m3N6pvWO4qKoQi4v0nvo9ArvszbhBrHrYKmpHAeOb/+s5
3jSRYyXMkUmb5xl4CHLVIFrsCZryfvobloOGAvnQLpTQUFRDPoHwOXMARLxKg+X/afJLIBpi+yvT
t0fT38y6qncVrJrzAnmon1yPWZK+uTpqJeUjfKVCMwQ0VnaNPXRwwpPQUqEsFxpoHz/+sYdJo17O
cX6PIZIFa25wzLxEgPapCBle/lheMU0ELyC0T5AFNvyZaXqlbWqUerUahLj53AB2YfAvMnTmdAIn
SOVvuIhAJ8TanUmQVKgCga/9RxJrrTIAadJGXYU3aO0sSaPzwkXAPsyFoLnN424JoaD/I0lzcgDy
zrrb87c5jWDEdTuWcS6uqVPW7ZK5L+SRS7w1lDVPpTMwJFnSZq/3f3LL0L+VXQJ8u6bN1H3g7TTu
6bAlj5eNzDO44qyhNSueN6EVR/6PIDiyu6Sh7J6LrzjJN2+cziZ50pOKTAJM/ZPNMwe0IHsIJTod
T34fEiitniH5su6H/Xm47snsno5ZZggIhj/dbMdEm5VWvDZM0jjCIVgmaudRCcj+uQqyjkOkc0U6
HP6AbVJgCv3SyGFuzLJ1fIxFQBZ8LIaFIX9Tis+7OY2iTrXvH7dU0PPgyDvxApumilVMBV9lnr+c
BpFvTZ2VriPRUcNOlxeBeL3YA100uuGgWuv1Po+vRzul3e+f3lnxCs2SbX4yJQ1r9L/ybvNpmhAU
bPD1i7FceTnJJ8VMv3Fz6Nk55L0ju9AuBQTL6R5Oj6bEvziFojlONFrDBDiw47LF9XnC/EwiUb4u
uUq0WR7uddiPIf1KRwzth1iB5YucuE+n5LUYQIFEnP3IH0+IeXUTCQcOGsUY3zBP2wziM9+6OXK+
8OlqyigyEn7hJxCPS52tHz0ix5yiP96ABpoQYubxKiaa+MyP5c9inb7lG4KxInIYRcdkhHO+NhH2
BpwvL9eldXeSa3WC8XkqP4a1gjurNYhr6YyiL+c0jb+n9JyaBmvcVKbxVrzTqOMP/NM3D2nl48Ek
4EOe45tD8WPECyScdXbNemRNwQkgWrWGv/XHsXjD93Vlb5+ppe90X7qHwh1JqrLHmbnxjZc5zqoi
9WIVwLtGEK/bWRIE33CzEXym8tihMbkORP7mZOsktCMzGLSr/1ACWkwIU2q9++sYQHYcou0zWpY5
CbFjLxDIWhKdljQSRsrSDPIIxkfPh4rLtpk0FwOrFTSwf2KAzBjFFgDxlYHhUmw25t+6AdxBWeEX
rvDpBJhjNeCO+3A1jW/6rnENLEesPeM7xNhDycr8DYISNr89j8JIpHHXrJkKkCvLpzepclZZoSGr
pDVU1pHGn9+Ow+miWqFBJM2TUc2DEPnV+1FAGIbqYI7ZZ7NOfwTfgDCCdfyuzOjYxrAfmCk7PHgG
MdEYz48Eo+WREKSlwvzRGu4Et9fuHK27ZaVp2PWcF73P+51bQH4KtaLjUJJAGt7G8XIgQRNiQ2WF
19c8tD7OpJ+oatKwvFt/z1RFwtUiBHlwOY8fkBJBTQ7urjHA9tAJHpObalORyhyZ4O95uF/bZKoE
2djO3zTjD+P1Yad9evhk3hINjhqo+qN7cSuX1dPPYr/KCU5lTBOVUCNVJo6gf2TawBGertuuh9Mk
cnR/4iv+xGoZRkyZmaQpwZECT7hCCDnsojaBPsj+dyQziXaEM8a5FvK448lZOjtXzfVMs0lrJhiQ
FjX8H2VubZXWtHz/aexwY5DFcj1zpNnNyiNBlNF2jf2RHEhjEUITpDi4bixE+UKU0oyqNJsY2VwT
Cn1bA7ILuHeUAU1Z8aR4tvLFyIlKpP0A4xlvGHfLcHnCWgD/99IO9DzQHr2Fw9pJzgfwAhibVdHj
T6zeT2kKzwuugQnrOI76TyqnhkhayUb0s3KtWE4cPFnspUoUBopCL7uJGTPjmxxBUmx/8GnXJbUW
CT0ThZxze/EZ7m/NZyj7C1vBh7kisO0QSanIUqafZbZgSKlR850d2A495KPujhspofYsSctVjrsE
c+HB8DK1W/oBuZEltBa2ClokpRzjJt/nAToz/BfJSYox2pXxLokoxFUHqz/0/e3Ku+HX75RKIK3Z
lV8ExCrjVeuxqlLdymT+klLjqCmuhRO4gAnaOeDh9cFaGK6rh4jy0x5IGSGmufyhzlqYPb1OqjLr
77Pdsdg37qQZgq9oIvvFGPpTw5WPUYK4XtetlY7IekG6Ezi8BIvBEWt5LO5+Abei72wjZJl/gKud
GOP2p6lcWHHYaAYXpVKskIQZWnVUBjg5JNvqX0TzWcZ/S3pa9ShIQ5ouAGLXRGRX23cAoQD596/S
RJsOjlqoJz8fHb+wYbIoKdLd9qJfqdNtmCu6Mc5Ct/9Upyf7cpd2tkO5Mc2Sq4ctt4Y7cMTghfbI
ZRNKvlSUT+WLD4/U5gx4MKOESknHAIvCgw47HJuFyv9R/CUgx7n3N09AXHPxylc4R89A1yl2LJ9Z
eVLDNFTcukoqYrXGdMtSaZwxIa85o+3u4ifP6lAnFIM6z8/AM/yxRkEj2R35hULoi5FXZbXFDBac
RaAuIbYzFx/WHK/kQp1f9zo2lVPDC1cXejv1mBlUd9hvwRWhPiQmFFSv219YF72RP8hje8un8vot
u4XiT9tnzs6ISWptSGan1YyZx4dHUjc9WxAU13RYuYQsgWfz5HnaZBupFoNaC8Fn6wXASXswxcdY
2/QPh8ZsdZKUh9rqeHIR7SVBf1lb1sOEBG6f8Ua3w0s6sy4VOOPhX6R4MwGltyxVF0BpCTpc6dX2
O9JKUQVMGLkrLpc5yoK5NWkm4qBcDpdYjysUTvXWrTrqeOxiYODUzvxbajQF6K0sIc7W7ymBUhPk
OSg5MV2Mqjp0E3awfM8lt/2cYv4kePjCGL3bAHKcgX+aVFQPF82ckdrQ5DIkZtieXP0+zQURiEgM
Sva5liwtBkmk3G9gI3HRQj5PLYv2DkcW6442gUE2f21MhQnWRT4xwnRPWWkm80uFMzqqIpNde6St
Q02Qnx+JES+/n9Wu8wEAoHG8wtyJVSeugKRMHU+/YFu8JLIUdwRv2AsA0XU4KAuaxrFwuL5UFCjE
aYvQPx1jyPtV2ibLeVW4+pHGLqHKGXEqWONcyBAUmNEzrsATh3R6AGeh8HTlHctqTiGgB0TDCHC7
FUqpym3vKAVBZKNo9j+tBIrSlpUV9jFcMbLVxNhARoSshn2GRco7zD9WVTTVqDOY8yWMQ6LTpkSO
g5QycfK+k68UTgw/k2uSpfbUmkdb/TUDVU0/7qL8yrT14kFGxbUuo2PlC0L/o4dS+J3pLUn293Vx
bqaWf9zxJcQD1racx8aBKggnWEuFVN4h412ZaiBKi3te5Kb1M1tgb1ncB14IC4xctPGigSecJvDY
qKquMZpxUq4G+LRJS8XaTW1vIp4vIkikDqdfVGI8A+0MtuMm0ipuAe69tZRT0AoW8gqwqTS/Uech
WPhOqQSe7p6PZEKfuemThY11LMXtiAFih5nVMzqeY0lMrUHXgueGtCsJhhnsXMU4q2plmEJoGHPn
w1wHvg/ZF15E8ghFniyDSzv1D8RWEAYouHzzHWKy32uWl0E6jluiDct+zhjb+xbC5s+Gqs+iW9z3
VNSoT5c+x2qJ3VOsGv85igMIVmpbiCWfkCbN1Qopfc6YnuTrpx0BQMYhCzB4EOJWEH2HPM0UU66G
dkI4xL8d2wTZnGXHlEh1DfmeqnIF32VIrHtqkPuHgnuBdnPK/w0aryYM9VzsXdOeMuPo85fAGeSd
2m2ZEWVbLP1hwEPafgrq+Nfj61js5dowb7sEz2TlTZfoWduWlIpv5BhnHYgzHIKA0RYufCIP8W3d
3rTHTumBqpTgWs6OqGY6tNABDk3dPvJVNEFpm6gwKiqlYLKlk6U/B61JiIukHdg6pHi4Ty05/Pz3
vXwuyFamWATdkiekbMY7lmY9qF8Rb88ssLSQVieuTvLxusuY8UL8B/RwxZkNCO+glQ6cj5ltxsPn
6GlR0vBNk6orGV4AltZZYX2HAGfIyQpGCq1hnqWaHMsBFY7ByZsPSmjAJzInMi0Kw0/RH6Niz2vt
iQMvY+umM3Wny3n2G+zTeQ8Q/NDVSSJaqz8nP9XDCjvdeqDPwe9oSW/1Ji448S/JszqwBo73yLW6
f++djm91zMr4VyDBg5rDtC2WU1BGtvAQIC+/fLHhHlKLA5t3KaXD/avT0MYaZw2jWX6ZaTxV5c52
Cb79/yx7MGuYBt7nFuKruiuRb53snCDq1Q191MpIPTErVwGdY0c/qs5eiFWosqiRzFLHY6uUKTEC
+bhTcX0I6O1kB/cmVVlcKQpUFrOQ2CSxBEHwm6km4OQ5pAGIKZWeDCe3fAbivAQEk29mUxI6D+kM
YN68kqvl4wPtijjtz9X7NhjAGkXhy37B4a5Eoj7129sLHjFhow7mZUVstgf0riKCy/xAfvOX3a6f
aCM8G5QOMLcfAYs3gIYmYWP5wVQQtVb3D3SISlk8XwSiodEF1okyuTYqgkaWR/j80dyukfwbHx1i
3s2JXa4F0L/SjkILfrfqpHsrLedd2DCNmoOz79MauwiJJJIKHUWZDQjwZWtwBOVre2YQwXAbdLEv
8AbxZi7eW0ABu4hMtapoS2VtgN0ZT5xCCnhYKBAQYYh8LNnmdvJ6XUlZZrAapHjFjU8wbuAPMr2L
ZPrmmI3V2LDwlDXUjcJ2nF6lGH/XPiDCvQf/M5FTGnfHJmjZ4VoQyHfBTKsj7uIt6WM8Wi5x9W0F
+Vpp2qymJeUEELggnd69LMuzA0kX0YAE3YcyKs1SYMYARrK3mSErvyJmU9e9bIOEfxF6xbDp234x
bRtBnIIQ8bMBsEJqO3TLyTxvAR+CT2YuTUbWuajodZcXgVqcEOz8bhbRH1QZES0xP1zYDlufZdZX
cl4Zq+fFI3y/EkHupH4dF8a6agaNqL2AM6BRuhQx8Ke1366ud6/1t7A49EOBFXMuLwJgIrcbv1Ci
oJOWlPgI/4vHdayRJ9l7zyFv1JwmAaCpd5nw79SuBEVHPHaPis985Uq2ikU+SQ4zudfofRS9OPlP
8pAZ8Dlmp8JNE4N2IEF0UCoDDRhdd7pkw0+MhUMtPHtnRsM+2W4DmxExHH0ND9Z2i1pFOwdA2tSV
HT52fo7F/EKmegUtf191kWHl7jnJfMRnKZ1DCY/L8mMfL8KWzz8nE3GLN9D/4wReQz0XOP5ejcAI
sHC3ZVjrw5BsdBJ/YbTAuOlviQmTuDM03t5TFtf8hE4K41yAMPc8mQkoIR4mJjLYs64miKmURvPV
y5vjTqlCgYR0UL0gTFbys0BxtfbDQHRbgEu8wtGW/sIfAT9s0jQsnW9AlyVDwFn9gBuwP1cUXMvU
R4paPZQBHvLS84aa+xaVBkeHCd5Bqlq2Rc+9TaAXMI9EbVi2/egQYN2vAY7G9NcXlcuglTYv6xXF
A6GBvVikSvSkqqxaXo2BAIjhhBBTnKLGE67fettt6O+xKr5WhSjoXfN6jFxaJ2ROfR8VBX6yT10g
TLtXwzKwi5mnDo/FfhTE6Z0HLo9VMNekybH4/cPuxNg9F8BrRH4ybFdX8kzB/Vb8J2Ku26SUuF4b
q/11ml/SysvQt3RH5Kfbpo9ygK85EjdVlvqF8BnX28MzQcOoCMbwNbcdCe5iYVBXr9HTFoDykaul
Y3tAxGE1dS9Fss5QFdoFCMejq9pyey4rbTcIJU2iBEQBpd2sFutvTCAG8pr5MlL3D3aqzYLDnXYa
8cekOMg3PF7J9thdS3ReI+9BQgefTq2+8Xf5t+aAiMTrmT852802Y9QvFvBXdk6d4r5Niout0VO9
nnGDx1cjW4Y8SxGzUu5tg/YwyWM++7IBzcHyN+PORR4jiC0bfnj18BZFmu96ZJzP8RV7iPJ5UHGB
shlVdDBHaJS/e9GE+2nI2kMQCk0GyC5gF4V6+1n7r9oYT325Bt07x8J9HQFVquP1J2hiKbrrNkgs
CpmsEtodpZ1DcJGOVimkWrOVpcNgD4Rqr5nGNyWk1h3ipeI6d3HdpQNLogJvWrYhRwC8f4u4niJX
LgmvZNpzpU68mr9pxL9+U0YK2aso+iiaRLK7hcYS1aBy412PdYAucAx7LfvFrkRnQIE8BspHq6ps
KaVnOqfA2o0E9rx/t8NJCz5+JUurSgX3/fTkj8hp8cpl9bMAxsEcVV77gEb1+kEW4Hg9OVK1a/No
NeiNapVJpXTGanlJkMyeTJs1qSM1Y2zuKPgTK73qlw81zcbzxucKDMMcIyBv+A7DynntsQN5SSwl
3335Sn1E7/A8Ci/qG4mq98SMJL3FL4OzWD2QoiqMktZWssrMeoH/pnKFLTv8nUnxyyA4KMJy/mW/
K/JxliZ770lPse0/Ac0ANleBpOnOg7mo6xRlN14z++R4TyDcsV1wbfTWLt6YFN8/xFCHdZB0XNmy
VS+/R5wOTnzskyqFOo3qzVDL8OzTnhtBzfjDUZS07oPXuthQIC9kyIfX4mP1wtAUAD7UICKv4mS2
xehWyHW1ClENQ9mXLTsiz6Ct2ogdr4KbGMu447FPW0sOyctvpDUwOIChPM2DAMWCODNrUnBkMFyV
PtROPLXZXkxaX1BjRv5qSPkmRq0kW59NOCM9DR3tMGKbscipwa+6bSi1DvK8xL0oGpAeV0FqNyNC
ZKTKmVjLSmca5+lJjFNcjwsLOmPntONd9blYSv4A3SMvPka/mhbucA5QPbWrk1cGJOOoyLmYZvDO
tDodULVnLnSbviz1ZWQteRadFDP9VGUwqokDnGlDrM1Wbt2Zx3q2UyBW6YIOOwN979DFDQqK/04d
LhySxcgjDeLhFJMpzS9p/lBh3V4//xNmFncqYM9qns/PeMfE1WLEL9a/wdPo3wz0oUUCrpOIPuf2
QNfQx7GskkG0YdQF0oiPM/NVXgdco2TA1sMJroT95qzjL8Knh0iDoe95p+ix79W8vnF5C7EmvumB
1f9AgUYwyOxNK0LfZVFFLrplr3uTGI+fDHZnWw5IqYoBaEv+kgP5RwRncPJPejqYCl7E52sOUX0Y
zxBU7obFdhUxgB7YpXVhTaXZG0Vtq7n/1j3xgUBp8d0Sft9Cj3DgO0dn7KWBS+OB7NK2kon3xuAo
iV+xUGvNnBdZd8YGi32WNqDk9TQQ517DvBurHCjqRxk2c+nu14RCe3tAbg8r3r3yTvTzjS3VivtU
2PJNSo4CWNPnv4IVmmAW3jU6X6nS8oo6rAPRb26lK2t8KMeGqTUWvFPI+7RSU3Y+CHur4nSWjAKd
ACazsE8+TLZmGHcW9KOjnRStzNL/mptLxDe0v2UVRRFvouR5ikiCa4OSNbD7ytFJ5RiyC/pmfus3
/Jtv2TsVRZL8TFolU8Zjb9MuBfoOu91vHp5TOIDyOfaQ4GiT6mcDkJUJUz45Adi8jsYfS4WXMt64
kre8SjH1SgMMxXNatkguVA8pEBbNZVqGaXtkSR7JG5H59pD9s6hCgj7CH0hjCjeh24TzUxFh4FAL
8i+a+Vl+08oykB3uDZ4KfgJJoeuSsTIzlN46ihCxOc62lIEmfqVKst8y4hd88DlyeF2T05+Hqoxt
LCQ22/5bXzau1fY9aA8owNbOfUNHt8vmtYoMJeb0uCrt5RI3rVNMDHt4QWXx2SbdVVK9gZYrnHsg
4O29kP5UvJb98tZF//5R/Ca0dGD6ym/G7Zn4GsVg2prcj8z4KqZr82in8rU8/2pj1ju0mU3WfSiQ
Xs3nXmau/KU7NUgTfKCUffR/+8FbtYC8ZsvBqCVCHSZQ6L5WSzOHVH/2fEVU4ASkwW6rSZmuAVkD
oI4R50/94Kk6H6oHnklVK+PkVFi6YMusulMzYtGcl9n76UC2zdNwSGioOLbBZD3jSNQGZKnd6ns7
gjEPnsB6aQfYSs2nLeBVXSWb3Awjou9uk9EIoppKpa9RQXZqtyGkDfN73tO9fVsyqqaoXm20lMmt
hOFnjmpUGALH9Hh1gjcNG9KluNceZS9N8VWA7193R2YDSqIWOCni9VdLgPpJsH/0QagVs0GKhT3D
4KDMN5OTp9vMsx0btHjTBZov69Z5AC/ujUOFfn578VsZGH6YtVysaO18B9toD2oaIGpPRNoCmBVV
vZoQUgzmI43n14xsnpIPaRjg7dY2Py5oj+3/XsvDvrrlcvNuv7xYgQ4TjhlqNEZWfekMTWnmNWf4
wd210uQPz2iOedd1N+5vnpdBdqFlCaxVFr6pLtksSJp6MFClKaE5vGYPweQvZfyVpS5jtfgpD7bp
3l5L8QaVt3rUh3O92RL2H1WrYDOuON4e8Sgghb60c6AlfgXcDpL6lir7PQLOwxFVIZ/iH8Iw9Man
X2R4rqiedHgAHzQssxoy0DSkCjOdobCESJHi7OoqGavepMRee3JMcJCwzpuatS74Q7lNIDJShiiF
2clmny/ngCZjiziKfcEhwBkJ6vV1FLjAHUvtbDkPXEtEgoq1j5bbvfaGO4F6y4S4ndEl8S0S3b6a
PJhxjsdjF/ex/EDPRzGiGWJdH0paOem8hPh06bqHMeHAvlTvvcon/ogaEFTcBYg6NHfgFmc9RbpJ
+31hbS1dxI/ji8W/06ujVuIwSKqOn40UilAvWc9OyHAfmAeO6yMLu3OVLPpH9OST4qNst6/rrMwo
Q2KaW2dE7zHKT5H1AfyJQxdejFRm8KDBH4o0UrmN8SwQceHybtDzX6lf5O1pcD1inwovyGLjzFEl
YkMMk7386MSNe/pI4qQUf2mM0ArmNxiB4bMQAkca9jXPt2Xo6gfAhrCcX1bmZ8Dm+Lv+ilov/bK9
A++B0h70LlB2Gi3FClAsM8JKXSdP6mbyFsKhAQXSvynj7rRzA0fTB20wzrnuz6nFIKn78X1mz39/
8oCjdTMRIMoQuke5b0vC++hVJcWqI+5uZA7TsrFMXGyEWis8KT+SJ4YKY8z4sO0J3lGiDyp3zK6f
gj+KVdDndhO7gpDgdWdJ9s9pz9yTxp4ee/VtGE6/hY+vVtgM8xdAokzNqb5aHoAX7SQ/uAadDA1S
fppknVJlI/m8oyEpIHqUi3ex0BSm0s5bjsfJU1u+RhKULhhaqKwKzFb7ML1jJs4cVuTGnk4JdIKa
40GjXhiwm7DgdzzT92MxydTZolTtfa6YfGfefvMzFSj5OaYRUDv+8MJg2kqJyvREYgup0MyQnjF8
8KLsVX6OOMOjBNk9/bLcVeGmjkxARbO4JD1pptTlidPaTrBiYg5uDK6CZVOsA1+KjEllh+VAPo8H
cXDV9J/ZX9TbOkfJNjV7avu5j60tKinnImOzFNBrlDJmt1eGrzbXOAj36ZPDbooWIrkqJxZd0bkl
/7Ep3jhaxDwbRmTnGS8bTE6LRHUv+r7f/itUBTGH8mpjUuqomxUnjjAUpGOmttZ0uwZZslP8y1j/
+HH6d4F2Y9pfsb6scnwau3EklmbULpbYfftkDpJcHUWMQk7A5PNr6Bnz0ADsdIAg2fZx5BrV+OqX
6yMZKHg/vyii1qmf5NSu+UROI8WNWBNc1eVfryIaAyf/WYU0LyVcVN5Nq6+CG5LfA28pblFPFniu
fzvm8i/GmSUjZ7xs2/vjj1Qij0FfLVFcMlDC8EiZLAJmGLucFam8UgKEUGRTRbxV0fYgl1SvIrf8
n3q65Zw5EWX/jPgEzYH4TBMPYbHD4/uFOvmPOOCeaAjXD4vcjaJ9dgLOYaTZuMppr0ZFDj6ZSNkC
I4J2PHcXTMiaTQeiNGGWfpk/nF61a/UqNdb/baZW7Y9YV+kDtM/dvcMhkmXRCyRGx3BTjqmhkkJh
ELgXVRLVNWaANYWufFbXqB88p3W7lEPEZTdtKJcE5kFsWsmmtvaV843RMxZxtkBeZvNdXkJmgSUF
5xa2FtgLH9A5NqsMyaecpMCke8pkS86aRofV5yt0JDtnLt6hJzMJBHFgYMVE0JnP0Ln9f65WQW6C
N4LxGQQSmF54FXkMuWBZ4L+0W2p11KGTJrhZbBAf4X1JoHcdW0jkkZkW+LnB3+vvhqZ26pp0nDuN
XdUZcx19AFDzAjVcoNJob/ok7dUuGWNGGZd0mDYq7u0srSC+dw2gTsYihEU0e0QM5LzSoHrnEAaA
OehxKuIRO8ic/dYbaBtSTWXGPbO48bwTkscWVzg/Au4TM3jH6yVfy0j5ds6CKCEKWZ35yC6tf87e
LhexaAFB2Z0QtYCs8g4Z7/25MbabYaO3kEJ5bvuWFN56w59giGrWHMm2DgehIBtvE50FGTgiHj4m
4VUBDbXfXca4IWyU0kddXlfgzxHKnn/Z9P07CS6MhNHK1T+nPlTqr0PbWBpD5pNTM/2qKURjSjQ8
Poa0/bFyuDDCARZs1qF9OPTPZtm+kwR4xUBo04vnZPb0PjFCIMmnAPXUgY2tnbUNkK6AvxkdfkNe
Xwq8HhtW5msXiUgME4rE7Zg1yUGWC46h9j5rKcLP/g5SBFtZFx4qqQGBb/pcs554+xCgNb1hW83z
DosPeBTUqnatS2PmFxoTC45JoQhujOm9y2QCt6lROd4LNWbs/b7qt59Rj81Rb1HAJN81N9OZq6d3
dWbM0sM1ldU3XoWF7Y6KGEVlVO6HbdyL7Pmb3uMKcWhKas4jqN4cPFwRC/JjR/zyUGHe6XVbXPb4
Ez8AsLFjNmFccE4g+3nWvBuVlr2cAZHLXSsRwfQW9NpVnHKBf0ZZrGwqTT5OvULWucTicn1Eruf5
cEqsUZ3vRucV7VsfZDbSmD5JyOSJ4yVzDev/KOS/I8KWeKTo/4KRtBbjtnXQ1XqWa+Iw+I+kwYeQ
0eYjjEvklXkMxi+www/5X9jdQcdaFKtgA9rm2wtNldi6rthjYfiNd/y7B3luNyfJzrB5wMB55+Wf
qPQhxL/jFB/MRpyMwhW4wC3XNjlbg6A3BnxKbOXwR4fN+6hvwc08noacJQUGQjfssHr6Uv1RtGpZ
TjGTE5zY+VnVVAV8p6rz1WLaEx9DwkOen66h7bUsvKnGr/Ng4WRUCUz+bKx9WSWIpGBfnJrlr4Rm
7c5sO59NQWE8U1BvB2GJUDhhfRQDOkEN+L+8l8nRCA+by4Nvcj0PdaaSs8FA2xP2AkPDQmNxorOY
CubRylw+lXHz2w11m0k4UZA+600zOETbTiCgO9IBbT/vaN2l6oYpXN8lpHLNkUGFz+V+8azGcKjk
6hJE1B96aGVlRGpFtoupT7OxgYvkZjhKya/Rpvl+MUO9FMtHbbf1GrnSeoat5iUG7Wbz3cDIjNeg
ffUK4yZcHeC53w24XtbCDrT4onb5/r2b6lP3TPQaPLPPC4NCtUrWS72liUegu1SyozWn0TWXDgGG
H8pt0xngQ+5MYJ1LhbbcMCVqCu5+2HJoVvQFSTeTWmjeKMI6UAm11V6D6DcBtPjU4yRN0X+6OWhE
H2J0n8d7bEOTFADBHBu74gPGHGNHuwZdBqwiyDmYvNAGo033QFrAOcv9hhg1VMTWMfhi63FBB7Ax
/gyUZW8Lne+cyKfA6EVdb/FNGXsfghqQELdGkKpvVggGUXRhbukw7ZTHzcSoloo70P5iQ3I7x89h
p1AujNAdSihQEpLrP6m54xaO0WYbX+LcsYd5Mnln4UONiVriG3wFlH3CQxJzXGMKGr6mAkU7nAKc
vOX0oE/zVBKnkcXMqG9S/iLZsdWNRp5V6HMjYANjp4VgaVT9d1MAOF7K5sGtCI4TEWVcPOxKw2fk
c5oaUYi3vGy3pmQQFGubjKvPFKOioyHYIdEZJZqd7qWueEzeO3OEtk368aErAZ8MOR7e2q7mXQ+H
jtooLX/vMNmZiSsRwGYI34eLhRsMtmWKPHDEXVJnld437H4RM2z93QyUh7JRnmRKwyqyLf+NFeKm
xtcGWs72WNkgxNyDuBbV1ARRK7dxzjaXTpBxUMcD936anjBXr7g21i1O7KkeBNiKPyKpiLJOcojF
uGjrZxgegOXJnipE3p+bqDK39VXap5YVqq7z20zvjJczMarxR0/7HPv81tRtDH218XI5XpnfMuOJ
NT6N1v7O+vQxYELM7tsBEXhoZppcWdjPHi4wH+wUcA/l5SrM2j+VmngfIYC2Mw2S2g2bu7P+SC4y
JeCKUZ46br0X8+a6LlrZI38o9HEoR9+X3QjVzZ0Mv8ErFrEjUZb3VvMj4m6GDZNax3L8sdPrUMVy
wWroDYmecjA6Aj1w9MqBQZhdUSSYKCR2MGMY6IuG3FiWdMZHrzc8Z8A6+Yue3dhdzi+43brAwq5Y
Pk9DZdMLy30hq1I7/24O78FdiXcpkUOT7wFIu5Ted9ajUOIO9wWnDIe3boUQzbspiRDSTZEv2IYm
lk5WonsqiEMyXv8uq8hxSQn0crcOwCXntGqcp8egIqCmXf7d3AU+8b8dxtrhl8pRxpVMi7SiPig4
gCRGCbKrsNaWmE07DHf/sPBTJSNd9XpJOb3lTPsbatbBmr6+e94YSSedeXLsDVwI4rXxJZ9eEcMl
Sxxz6GToswzfLRlX6aPaDQdnFbgH8yl4HmsKo80uO7FqUV/wIjfws41qxyoCET2+VQaJ7wUuYOu0
meLp/e0nY3JR2NCOlpOJsXH0Xsc2jEELVBoJ+vacvS23njkboCzOTZAJMiMUPWnr/wfhDXPLrLCM
jlhr65LAz9SnuO1bOo+HFgNuOJ7unH26nz6nCwE0Ryg1wGvZ92bIBC2h1Ryn/WDOafvRGbtCSY24
gOdPjuU19FC2r6ECqZ0qwklTJFILgijhpnhuFNUuM+fNAN9xsj3Ewx4az3DZHUEQPx2ezRpZXV2a
n3sRcw+sWprzg1WzFclKrbOB6ezrhAzx/2r5pEJqBlLYWkAhipPMz1MPRWzkEDm/IKHu3O9sa0/Q
WsCOn1jr4eb8irb0RfR7SUcXEYPwsW6Q22u6Ow5h9w9A9kYNeDtu5SxSnpoWHqCRL+gULekTGs+y
97WUPPBBraaQ+Jf0M2feo+9T85xc5aMt+GRjl0ZNifU9UDVAmVN0P2lnbzvVLbX5fmTfxd3K2Vd2
byeq/4gKp4AZXIITZivY2IOcejNTXVBe6OgTPmFyTQQnVh1eYv00QB2DirATa58e18DhNZ9aqnnZ
X3JYLV4UE0w6/78SwBKvotNxi7sUWzYezNgcFxYT9wYBFDnC9NS/F+Eo8s6wZkuDDOp4ewBPXPeK
MPK6G8bZrOyqWH3uTF4DqMKjGcVFANzZ5vkdLo97wmaBbhgPsC3XpYqATRkRkplZOPBkGf9hcz02
Pp7mW27xBcy+lySDokQBi6LhTm/lnpyuEPN9P7aKyiBYoW+BR7QlbfbrAouUPu5rlYFq2WK9jZVT
CiFyvCJwvDwEBIABHsYup+QNSQre0YMhr/i2n7ZRyGvJvVygf7tJmf453cOCVeIlY7quoHXzVTCW
PTBLd2U64HN1586yOOA/8xwGnDhefIvaIvwHPVIwlI6U7Q/olqVpaXfp2T23iQy1Qn6ysEJ1nb+c
rTWlCqtTZD8lQeImw2w+u+o9b2+zheKUcMkyKfN43YVaFGnbR1X9ewAJky7ltmqWPra5GIP4F08s
W6/nrejV50XFtHyW2CtBb2Z5fhfJKU/XTJ0CHgoBmk4wyvh0Sq3ZJojAwT/gzJ2D51HXks/Z1D9+
feoHPmDk6LfXlSCVB/Abnh+HiuksYyAyFAtzj0bAtWuiw04uv6Pruc4Gh5QBxDo2weCxsuM7M/Id
79MVdJnUwBI/9DjLAWv4zraTvE1ZbWENyT7ewCJmlMFA1ea5wyH7Fj/t6oHuYS11GBpRDgSN0nHH
c3r2C1RI4J0ty101PhdsmPhzA0TYYaom+T1t0uJfmYgyQUTANfNDrUZVbCxnInlvKWcxR7jmCjS9
isbd+Z2vhKS2p6k3ip3fQaTdc2aPY7BN/K+XfGcZhkEx3zw5vG63Vr98k1v7rO6xLvzhHFG4WDiV
aQjHqzA+vOOoxhHugDii9PGz06Y5R0f4mFAUO+4zvfefrFtPn6AmRtUz90YFTz6HjoSxkilE/PNS
A+qXzPtRA5TnHeVxAHhVtwKp5I9WeEjpeLq+1505ED1ZztSl13rAsYTmq29WqUDlyAN1DwP7pmzt
4/oHw1xYgSelhbeiYNa6T+KnLLObhrKn2+M+8c6ygPCnfW0jfS+MwQ6eHijy2FZIpBcFjxz9ut41
gWos0DC892TZT8m6IMxzdPnrePhdezz45JIVsxMkSroe1m8f1Ae+7Km/6GhoAeXpQPxHFLZLdxvE
bRcolcxgqCU7EGj/rino6WeMY/zQZRvPP/5mPgA38LbqWeP+5pJjrkk2PzYST6UY/APFssnzabJZ
7GNK3lkIoJ2W3Tu0tcrT1SCmaABnwxlbVd+e8EANukEiorN3q9RgV023J7hNt8hIPQ5+oO47aD5I
S/upZ2qOGKAXHJLbx93CXDXWAvpDLAl/DV+ZWLBjacBoU5EB0/8eXeb4HNmN40xkseC/5BAAGxlj
BfVD58vEyu3GO0sgtaMG6Ec7mEFISa/rvInzyDRHyPo8B2KmSVZgUvcy+El7X/+caC8zoRXoICZx
M9ud7Hcl2asuPxOiR0CIS71YbYUysDj5SASR3atxLvNnm8zhRejPGOu7YrvmViHr98SuYoittIRd
IoNuqZTBBlBGgrZtjN8j6AxVi87e6UrDP++Qtn4I6HLVXkvlopn4RPz+vy9D/bx+Khai3RptJL5B
B2q0M1GsmBM/18y/eQBFTIp/L7PVvJ0NEkdqhjf3E0f4MtkgE/pi0eNda14La4yjNgCn4Honk/qf
i3324nucgDuH1/awAFz3R9b+S0qadexePkuf/hp0QebuqXhEKfcxF9cGgbzARYAlMT0kMAiD94Hf
W6s9pz8PF6m9d1ugrgpUo78AufYPHfXQCT14tJXX2JpHFchVl5hTU4X+n1Axk6jOdOrS3GXz1wsX
QJXzE5UyGhXDDUFjgKC+DK7ST+IPDXHJVj9sJdgyGwFm82W00JyeVnjgUeetlM10I1Ysa+UxAk5+
5aw/CdiPc8o2Aeq5oHMP9ptg8iUFuSKbi6m04T6dI9PnDUzsTHikN0AZtiP/++yd2aS2G8f+9bbJ
/o8A8DunCicpYXH2VZcPtv7t9NS40FXIjHc6deii3wY2xZrMjoWYLcidG++4NfV1hL6g5Jkc9spL
69fT3zaakEH/mlYNuhyzyL/dcKNwSjCVxx6QwFz3yUEG8hjGn2CeY4UbLfKLw8mBYmH0QHi3bYvM
3HawLheGOpT+2dKB9ZO6DBA9M0r3jrgZU2mEoyQXHhc+C5NBT7oqegkWPBnBim6pGtHzknqyFXOg
SonBZUeMNbWJQc2gZAC8OmosVxcD7nKcxKzWxEqLo7/z3h4QHkOTbqThdDXxv5ANu06Q8MgTrbmH
60dXhVP8Nb0zWrZ5jN51H2MUxJINvHBYGWAmzf3ub87fA2Se+n+gOl3GZxkXNSb/DFzxI5US5G8y
QQ9oUaCaAB18cUB/8xsM6ksytRUMhvq7exoW3dZclnCQi1kQ32dxBbeMcK7xqgacA3OagSp/71wb
C+N4zgnKQSg3MLBw3CeRBXifI/jL0HXrH1q1jP3XG9Xh8JuRoNu37cv8H0Ui9BwUU+X+t4G/hchw
3YOoouwOZphh4CjdTkY07aAla4jTnMupS6qKkQrku/ew1qC3D6LJFl/Afx5To1/eI5MBj5Ek+aOD
mDeW3jWrmcmDNmO2Xgwpn6wp6fnZErptxNg+qrFwnh392YAxEDhAU2xXmyVIAMLoeoUoksysKpS3
8yuHOkr0ZvrfPzDZzacy/nHB11QBgMwdM6M2FNYp+8VrX2+gJpOZgSwjX1o91yZPawVRmea3BVDP
LqtzYZiq15Mgk8NsxhP7cDlSO/GVbydeBGQEIj2E5pjpJi8eLlla7bYj4X7ZcMvjXPf4AG4DdFwz
cz+MXFJmtcRJ02VlpDAyn/93PWiXmi+S5efQXo4oSeRW+NNyn6TUTBx2uHicFwYQtZ8h2k8z6MCw
Jc+MmyPhfQz4prsblPFVW/y+L82Fk+296NF/e7NOWr3ksDpQzOLO5PgUf39zwPgyMb6lfHP1C4Ky
bm3+IQDjdzOc0d68cSxFVL1hBZpsB8A3tiUi7SvapUkG3cTmZGSBNPt0pq6J7qrcWd0H0fyiiCOc
lBQCPF3DRBGBCUQnYqnhedBw5HYfd85TP2fHsPzZvoCM1qSoUNjZktAiUUL0j+kfiN1vZR5vvIaI
vIyg3qblnsjpuoyk0wwArEmGiAZaNwTFjp0fwmaFi6gcqLv22duxhK150LSnin60F7LyvGiU7mWx
iKuG+XxTmVBuIWrlmIHeypDpGfRGz/vcpR80YdBimYBBb2cxQ4q3frG8BMCdmo1dnhJjVIDIO153
vykSkQLeN0CRePAT1Ly4kLVF+Xbx9o1QAncC0yHBRQWHn3bYhnuRJkcl2FvXN9kj0ZNLzJ+OCj3n
aUxvSPEwwRcqPKY5cFeeNdl9kZrSxNJglAlkNRhsG8FyEJsW5doVQxud8gyOjWHjLOR1yIfkB+Am
oCDEuLurnblghK0BENblJh28SpcVkGsjD3dPXp+RJu/gt5tL3PB23LAIcNz223aFzvGMqxMQhIJs
uYkjjVR2CDg5mxmeHsZYcXWD9knP0SDtYcD4wPJqF8HmvTFCZBDVo6iazREjeNUam7dtKUj5vYyd
gIGWrxxUh2hCDwENUBlxsYvPLbt+hW/Zrg72YTMCDuavvVxUwMF1LWsoc8uXvrSkB9DD3YBdDCv8
tf34EAul2Eqz1sbORiDoBN3zfACaOKu4UwA/JFldqG0G85ErxTm2KPxdtPMHuErQp7i1C6SjYHCa
LgLfmXHV5RZiZ645Gy6O/OpdVGj8ZCQa0HEDPuxeMBBmknFmdIwez6xhe/I9opXxcUIHKTNCyVUE
trI9yiio57CekYS+UTyAWd+iaO4z7wz3nsKMdPtW40Hq3CpPED53kcIetmcBKktSzu8k4FuY6wC/
WQ7vNfMyjZ6Dbjq5taKKz0gYOMgJ2thLBUTXnSUNtO+0LXryFlTb0+TrhlIepi/dR3YM5BoOmr4F
e2awOAHC+SJavthhomZNGSeFyuyZaX96f82ZwCRpNBtIrl/HIsmZWJGXLPnrXPx3YCdKQV5W15xn
9f9WL72f9bvCwKCxo975JGgZE6eGPSNJDPvseBSulvAc27nXT9c7SxpY4qKD2HnOgclxOl0ZkBwT
ofbeKLDxNnoaOnmJSn01qV+92ouDHAmud8mV/lsvnttjoJgRvDGSOAzLzD8Q8VuOmR62RGBA3OTu
RV83kEEqbs4wK0Gxyih1k4zO8D47XymExC0hNyiI9ieREte2AqgOt+5zc30DUkz7rJzGZ02VZxAb
32QW0ppQ9CkfCazXgWHd9KOeRh+MJsDld+a3893qnugEG+U+9QiQ7IfgDEkg2P/FkUopBNiIxJix
3p4QFpShoXbYKwfFU1wfa0n6vB9uL6x0UnhV7U4gm6ZQy9Tv2WJnQI+yXJFu98qOG9oUphJgZa+D
Lf6yFiotISR3eyorAzTPLfYNtdZ6Eacmci/2H5XzZzSzvJuSmEKJQohcJVH2oDBRV95Y4ihnR7oh
Ij77f0j2xyY7F0+b2RaMA/oYFcUCGLYNHxKM/1+8oUR8PKc+rq/+XefnYDm01HWGOIuU96HVcstn
dU/sd/mVDAjYptU+p8IOuhFyLHIZ4bkOtMGTE7mdkxXUF02IRXvvY+WBsZOd+Yy/zG+wxof01Ymx
TOaCtF3hcLOWI2jDOttL6DHm4QbyKxihNA/oQd1i/uV/iZHIWxFs4/qlWPeX+Ww2XftNkZcTS5wN
y3rjZzxm93Fx8R07gQhe3qR2sTEAD3r6zf0i3P1k3YBAfay0IXs2p0pAL4CvqkmNoBSw1UGCqi2u
iet5lV93OYfvcGUgspdO4HgQtlc/GfNG0BqaP7KNS5PSSZDvGNQE5BArTWIts/xw3iYu4SqeCleb
qrrpRL0DJd7TMq3RuVQVgiv6CG3bzBgsa+tlQuypE39fluSDJ4h0tUCyFq/iXQww/R+TGtS1Myfy
98xXstjhcF/5fKXeDgTC6fZMub7RWW5YvYhkUo4E9sPGBBl4uuaOyi4gw239XhyBrLghqpLxjiht
emyzxwHAQ2NF5XyWxbgIXsfIAf/5beqBkdxT5hXaNbVUx4PXDn3tK9WHFsDMb/eudXdiBoI0W+ua
s7xmZKda9cc3X3KoJTes+EDfIfgK7RPeTdhhSslQSbEEdlUfgWT0O7ZC5VdKrmIz/M1lm6tnIuZB
Pw3nhPuPTTVjxVu6DHSmBDzjYNrRlqiYqHUrqVYKrHHdrmFVjLGk5F4WkLlSQo4P5ohViBFxxk/I
QrfU56/Hr5KtkYWGImJUQIjgz1tmzGgACE9+O2ZBAmxOn5nY7XMagXktxM8sdzD2m4hLRI3adMGq
/ALFX/0ivayA185dZXOuC6+jAqPxImgsi9pTL5BpSVsnEwNY/A61RslFowBTHFz0SHF6Do+tDk+2
uWHQG9skVTgu49A8dVtBgRfTQz5JxD77W8B5yAGICkUjpRl+wSK6uKep9uWq73zfdF1oA6rGuXsu
SO/v5i/VJsltZ6+k15rdgYlRgRzs3N/6ciQbZAtscIb7EYlD1Ol0E7S/aJMJti26eDBqibeeISRy
HuetqxrnEPYr81D6y35XU4LJcPu08F25VAXBV0Ih+xh9ZzKpKoCb3q1YW5xpmn2KGejWYh+Mzv9O
CAPuc6tuzryimfdO6px/m0SOCUsiobPbnktO/+ATLpT4sGeD43mdbvfcDCd0RYMPNkGqDI6dGYGR
DRSLW5SZt1zObkcljZJjXKaf/+kdXm3gbC6jtqZh3kA4tsTC/xjyttpaCJj3u6NikXeT5lSm727d
SxMLWelYT47mqR90CrFJc1WX8vuIo4axGcZJDxlFLMn9EEepmbQn24n3rqm+Kf0MVVD7Bs1FE6TE
Ni+WmzS4/HV0RyQT8sonQi/2eNqjFmUBfZ9tgu7+a6rQg/cNs1JvXx0veMX8FwBjHIS6/lSqazbt
IUtdNbLXyqa695hi31nppkb5gC2fltjod75gZNQ9Ujx0OOy3U1lnrIdY806eHHbAXWCRxwk4pgrs
2YrwAf0dQqGwUlUE7frCbnNjyCVX3BnpPpuxk08LDarQyui0gUkM7uexCpCtoTgW2EKerSYVB6lJ
yRmeF8/ZPbHzx4qwpXpYSkk13TzVnKl9Yzu6x0zTW5MkT2CC/hMGRoE5gNJagpySxuymOBZpZiAt
k/DqPdQNxzlvUY2V9VL8xQx+fLvUAxMT8Ca6lXtbGJfdvPpzJRSq55Und9pJ51qF47lLVtqWn7Dv
YNqfubWD7P04ElROUXpLUHLarwgxGEvE25bS7bxYaP5oiJ+l794KzAgKPrwXJqHGhUfd6UpAKnbu
KK9bmEdmnj+zh4vBvIBO/S2Kn/tQFkoJaJNKG9Guq/D7qw6OK/S9ube4FpJJYF7GfYyLIIxIBq7F
EmETlAA419Bv/RYshBjNF83/x1modD5ZrN8/+o5css92LSoqA9mLU3A1z6mmPNvS2WWsbktwHMsf
4AXP7KCR7iFZcmBPTO3oYZsfoq+6EKMNfi09cshujCC+cVXeVOnoor2mcUiArMjTdr1Ozb1ZPw5k
1ctCa0YzgqzZ70fCmPQepsshqocd5Xe8recSfyGLOWUbvo/xitmY1FOOPgIeE4JVN+3CifoUtzhn
72Sq7cUIbAtp6Ff+DNjkLw3GBRCHd1C54Y+jxmO7yx1QkdWbSAakyCtOZTOIkgNH9tcKSzbmncrn
GD8bBl27voj8LW0Nqi/7Q+dF4OGGM+gd/kFHJfuq2/N7IQdXtc8NHcKKNE0r515zk3pvY2Vb/c/n
jTYUtKKeWnKjeMFFufQlfh3halu1Vv07rGL/OKKFyvVCqymZ7p6ADf6hHmrH96Zu9P9Fi0wKYT1r
yNRNJXOj7DiZLj2Gd3xWhm+Z3TUKTnPjHfuLWeHfnQ5p5n3VKyOJHDUvCtXxHgoPpXIzmJGb6aLK
I9CMy0Mm/knEPLo01tIDPAYsAaUEsgbGQ8/v/+hLJhRGIl3zFm7smvPVzfu6HRqbNDHr+A5QG4ef
m5uTq1rakAf3vm+guT4wWDIG26euG019SvE/msqC3xI9Rfzxn0+TDUM6lpMjlDk1hmQXOHoi4JPG
kbU8f0Qj1Yq8V1uPgoRMYnfIXulrTpLehe3c0Ben9dB1AHccIMj/BA6xoHFTcgowHq7aCBBBjabF
XQNPZev5ygxPoyib7S05jnrKjGsTFvCA9ZUfBPEs+ygXumFph8NqxnnLj+CWhY7IWMdW0tt7KLMh
JJwHRNgefQVA0ydYagfPe+g+0GauSV9HocAKanWL91wMYGxBWs0kfXHYZmYVCvOWREfhnC+1ag5K
jzkWl9PgUBFC8B1eG7jI+wy/dnybFex79/7RwNoornBsgRzgMR4fDCips2O82CB1zZhvvp4ISall
muL4LbmqLrQHR5wc+BmBGUuxi88usLZIJOhS+QzbNxbjFs8AZd4U/brKk9g8R5vJOg8UCLJIon50
zmWx2OWfEPe39WS7eT/BTTSWdYkau0ht7Uz77vjh2N/nfIhimc4+ByKXkes3PcCv5U6ZONtfEbHY
EQqNhBjn4N9mbCLst5TCX8HBNGezEmWl9kkz2u8MwGkoJRKUBTSOmy8rvPPMzlO0ekHIudcwh8j/
RAp2H03z3WTCifUgLj3S2X0+Qtlye9UMmWA1UrA/QlEchVL47Su5p7Jt+V8B0C/RChLF8SUjXFaC
hvV3iuR8KrDyGxGhBv/ZdHusX6grHKtFAV8A4rE4L6UlHiQ/CI8DI7qkOyys/508wZzIrz6FXhMl
nO+tmwHE9+zFdRmGctF/LUyWdSzPTWgC1fNlJcU+49iXxm7P4pLlraylPSwbvJJT655kwG/A7TTk
hJYtav5NjpAgxAfVW730pLwFlzv5z6jW248GSrzzNi7mWhK5yEV7PsyLm9UubNvNJTcveCFNLuCF
EGJUcee86Ee+EOLlKr5ntdUGUzMAod1MVYT7F/nMA3NOYtXLWeR0NaewBo81js1RKPDA7mYmjK4q
16jKKbykssQarbPBBCXoa4lJ8y0yWYRYJqs4ATU8nGZTitt464ClV02ANFbQdwgR3dM6gqbOMyWz
P+zPLNZQZ584EwCcR5af4ng/USyT9yMMi7H/jVctohDF6kyQf0IBgbLg/W6UawK4gUp+Dwpdinr1
2+qr1t5IaDHmBvYCnkzNMbVa08J5BQ9mYppypq2uL9yWfjtWf6LmfORGN8tDKTrgsyr3a232SOdA
imQiFpwossL9j94pds9XRIlRgvn0JcuJsVKH38DLIhuttD62JB+h9MrwAdcq5uXFyEPHwljFA8tK
q2yRq3+1uMSQSC5cCHNbgr7K6kgDkBO3AMP6L6wQZYf8l2NYwDvaNjNwDkWETp1rW23FftcjtDsi
bbR9XnuFi4gLTBiWQ82U8RDH6MDHSL6D0r5OUBZFRuDfvsfjazdQVq8OVZ+8sKH6pvAlBX6WZM9q
YNgOS09DJkUD4rB+f+tjwk4KuNyQ88YnbBrQlemZ7ujLvBE2Nh6KDgafwPhlpYT0XQlSf3EOQrLf
b1LvAJ9QBwST+ZPlTapbtLHq5gHi6aRvvhihMiZha29sQ7tBhUiOpUZYzyQSHi4QWyiLor17b5qk
ACAs4wlU9mWmqQe3k0PSZlRVD33Tt4/Yy1tjeWkFENw2mf8My0I1nQ8Y9CQswoN1YNgEULyH9Oot
El1vtuG5P0z/oBb9BI762Bvv3ibYKgh7azFWQc2Y71QNITRMXfy0k8KkqcX2lPi+KTbKzOpej+sW
XSShIS73hfju7/TW/d7k3lp2P/PpcMWqa88o9c5KjO6XiIN3yHys+jc3aZNEaeGD3TreCAfJFmhv
Dt8sVL+Dj05vE6B5ozgmEaQYxz/KFkeHjyNZyze7CqiVf/HXzCX70cZ27byxdG712dYU9k7UtFai
/IuE/m4lZiAjXAoUNJyr64Mr1sQrAAdvm83ftuzqLWXco05H9LdYJlI9mHOGpr9fU/QwSbJ6d6g3
NOZlUVkhFTiGWfM16cYVrvQt6lXdMSUE3BLawDfzI/yicOqs8Luhb2S4C6F6DABW64agXyqHXFJv
o8z9maW6EIhxjsbxTgctdQXtLR0JdHcTU52O1nn1kDPs1DIOTwR/x47P0Xt3VrViBtaDsDSVm3q9
zw4uBQ6+TDFgOjq835g77yZA15/gvTQsYSsGPbdrxYfl5hZENpG9brpuZHgzHN1++U7Xqux1o0Zx
B00as0g78pDCN3+FimxTa2Ny8ZUdwOVUnsaGrksubVKJhmSor1uI9OgVQIbuNolxyeVt6TR37M4q
/hiiOVylRXSEmoBSV3zuxin3El4fAZKnM38cAf7BKbdNxIbhvwuhgAlEX+bMIId0scOdx6vh/cgy
oAjtqF2R6h/y4n+pTCE+g05UCub79n+yzwshd98WwiWbtHy5e/gz36+PgO7irAHlixr+dMhVEyUT
khN3GcmybRxuYIgNlGBcEHMczRLFI1M994tMxE6ihF2cYmD1TaVHOJ3DhICmWianMJbTXtJRrYhi
ll53K5EzxeJVz4sJOS6OlJBh/xkupi6MIzPpzH4SddQC5Xddz38fob7bk0d0q/pVaRR85lnoP2MN
pv3x/JuHKNxVgNHncoBWLuWtlLz8kXK5rlLr5BjVyDF10+PxBpQcm6kqxextaDUwB3I4Rklm6ARc
davgigUR/r9zjxSjLz7RXOdZX6EvDQMVqoU0xMvfaX4EtpHRVZ1VoBYdjSr/FjX/AFMw/5VkjO0n
MDjPq0RZMzjzfbjgZi3nycuUxQ55/nVyGjUsOw2JiqSXghY7RZvScyQOs6GzdeSn9Xuv380Dj3pF
woRZZeCsTztppgMl56UPSY0RbszGSiQq+J8BU1EkaHEG0e4JZ7ll9H7e1kpFkmQCiyonf34Gtfc/
RDgXpFJtBign7lhbqmogeXKIbrb9TrspOyvHP0Gq+/3zdjrpLltj79mXCM8ygeH7obPnsMRjSRy4
vMRLkZoc+FTnr4S5mP+UnHQ2/vzKZiP6GFeaKOwWOcHifzr/kiaQAVd5goW2RjSwqAq8R+CDosAT
b1fjif0NoNH3QWadjQHsDpdE7VpnOxcfLdO1YckmatAT9MD07fNzAEbdH98LEvwqzuIEuYhNDien
oDkBRKJbysnRXEreqa+NYWHgUE/jdqQt4qh4HUulUwHexWxxrVvp8EItpbKAGCZa8fGN+kVL/NLQ
X92PjVQJpjk54DmWJOwP1CP2+bMFXFGWE51fJ4apW38VC9wvO6NClUJXH12qZsJG7baWPEUN9bSd
qUVPt9c1LUzxI5A8sICmskRlGJ/yCUt9nbhrTc7QvtV2f4HHQw0Whegi4CI87wYCGKPALhb/9di9
xSS+PYlrXis3yuD7zrQKaqFJy7EK8ITXXnywD3BFK2fVzNB1cLvWe9iJijSizcfksaEIW6+Iv5KL
AK+BJM1ExViRO+uFEbqBgB6y2KQJZYeTsOwN9ZPDwCOp3HFXsv/TMKKaF9eDX/mJXf13bsmkfo0D
TVSWQkXnHe0mf1Lfo23LuZOH7aRnTwKvI/jE1Dw2wcXzKC+FxfWyqPWaGFM58cw2WiStX6yvgAOd
M2MHlSSwDn2WsoShRh9Ub8K6Bku4ePzptUWd/50DXa9o32/ezB6ckQw1u4shW1k0GrTpBT183bu1
PbZfcUeEQ4QES6zQepmJiKsHcYUychYt8aIAX/GgwPrVfcdj06pVxTzBdfPI/M1rAed4x7GeR0C0
TBKr507G9LtqIrOX010u20E2QRPv7hNnu56IA5K7Q9PhJdG5v4Z1cLpl4hH/ZkeOwZa1rSTKoC11
GyD9kFuGP+71rjd+cz2MbjyPHsfTPXRB+adXJpW5XOImQmm/300DaWj+wR3IqDM/Ga1oYnioscrA
dIEp+G0bZlpKDBymrP9QHZjEzSukRNQ/bq+QQLO0YTzv3hS3ice0x3cLo95mmrs1tt1cZOLfBiA3
i0VBzTNTgLxFXPauUaAomndRaThqsZLH/tegHdHvVvTVo8lKocl+OSm49uyYJFWaxOWxs5a8ZER2
8MhxuoFHnxNl04UYSQcr2N2pm/9skiK9yRraKNxD0tE8VjvPoG2NY4Xpccxd2/NyxsC/WKilryfc
o2u9fPNl/6XJQHn7ctlzQjgC0G/5thHK0I6VzZbQUUytCTSuCKtEWT5SdvvlfnyUcfrwZUafTBE6
ylnY0qwkKN3Wx+th7805EBc0IwD3Ru3atUhZ+L4G0G37ndzSAiqGde0KvhSCuyy03AtYHOca9jRC
rUM+TrHcShG8UUvVP1x3kae7SAJGGuUVp2+GIRP6uH1sQbAH81loCb8JpOKGmKOJ25rGhEizYLbr
xUOKnfsix2EQW28EVzLw/sDcJAgcVUGUSKtpb34KgIU7p5Ndoi/bO065+Ny3sczEC1LNDDvxe8H1
ZNP3Y3h+VYuE22UFmlKJk1qFsWdWxO9s7Jy0PPePEFQ8tJ2MB/EPruITcuXM6G4qw78mUjrAkHEk
osxTBeDjaTLgBgChWoG0AvDVK8I6wYeEEsCrp6SrwqeJQIP2J0ZD5GXizthLbG893VXys0bvXkc6
TEXbSBRlMcn+VT02uadsomGZkYaHs0FOqGA96UiqATxc3oXh4THYy5+ORxIooGLox5QdSJh8GTkF
slN9fJvDNOt1GPS4/z9AZqNnL27oShU1w3YPdxKu2yTnf5b+fwb/nU1ald7T/jIsA4Lv8zyHZqxq
ttgzRcvwmQDzswrlnPXIHQUNOwJJ9hxo4LSJ5iBbRJUFDFKhM7YYB+4CvrN2YZJ09PDdafKhJwt1
HD61MCTpf1PlrENHRzV06W/ISttZ2WxCe+DQfXRGo+nlt+KB1TT5trTPfxyRxqEBGyRVLU6Hnn9b
N5PbcW89cvOAdZpEGhihOG+ftg667t5lXkJsF+gXvsW0mvlnV0V8iuvYPM7j23l8W9auAZygDknU
vrEVJGsxShqNXsFHaBXmBLC5qX4zi7d4W1L06uYzsGSpaf6TWDbaDrnSYOipjxwobIxPUYOczitW
YCesSWZood3Zv8kwWWwQffrpSygpY42TSmApDNexqvCcpSA+8WArxZCMai+FXR8LwwSv7ezjOEDx
vx1Pc/NAAqPgH/OXn7cD6kRAbiDG3RCHzuie7VuD9W2i8ESaM/hhEoLRf6J0y9fZif+9ud/Ycswg
+Vf91HeQ8vjL8+gzqCe3UZcKch3XALNvWwVnHItNfb1OR9fmjpEdErtoEl3sp7z8YH8uJMDz7WBF
Sf/PZ/1VbRASQuMsGdLxkH4dWCnUWRADBEPzNCAO/niky+H7WJ17EayXmGJURnrOob2MtMQrTj84
3TfIfXSa6oJJgKtpDXhVxLNFhvMvH7w222eC+tFFILk3PD0clO1o2maiPUonWGupJJ4dufxS4yqW
gfzOEqeQ2tQf77Iq8uWQlX4MSE9lTUkLQFCWcdGU8LwNRW4LYOJM3kmfmXLTWhV7JsEU2M59tFXF
ZQxOB5+/zsB/fpUwyztk7X90xTTVgk2esmEM/qkzmpZaTXEEOVN0NosaKhYd6BbO9d8skA4HGf56
Oc9W9mu2/CbWLNVkB/ErYGKMGjIyulVD0AJy5wiaiq8EsCfNPdUIwEOvHAWjPuazIpk7KaEOkBik
0y9knolznSE8jfC0holtHCQ1pd1oFcXZ6HbqGRY9rHOO6xxqpmXJ4LpA68wKOsb0lzwukwXhd08r
22AQ166FVV3E0VFqMBSbAEkBqKY/ofuzreVPTO1DKpvae7YPFDCzEPaa9iC+aSyKo4cv/fFMZZHg
hcOKXn8cTtt1lNvcBGFVd3SjxJtC7fSj3BjQAXrt2/fCGIOVSEgcafMryCu92aGFdkwkJkdvcDbp
5S6m9N97bFadDHTsQPx7Sm39Gpq+KY7YKhxskzel75R2HUYonHxRY8Fa6L93LdYGLleirJKnHILz
fjZFZLrLpIVFzhWzT+X/rI5QitmOB9wgFGST6PQcJ1xWf4yPRcv42sPX0dnBLJ/H0LTXrHIwsRMF
Pi8AEio6A4ykcur/Fg1ZXn4450h3CRqQgO+DiT31k43aB+9SXFyqYLsm4BXYb33OzjZqzVsOr80X
q+8V52U5lwbJvBQHFyfiQEt5q2d/B3vk0K22PFEt5s7ZXMu1r8iWBmDCaun5RjPVDuFgn43/UfFt
bcSIbrk9Qujpbx+Ma91RUqX6dK9uC9O6Bd/rRNKZ9JiDzz4PwmB8tuUbE1me6S7ROFSqOA3IIP1c
allfgLb6gUKYDNeFHTCbOVutEXMxiRc1Yz1U8hTR62HKlfs3Ws8ZZbMwDrOWANzIIdDA7M6R/Bm6
B8TQs2TMdSZHdqVq3aLGyhaGwObebkiCzC2PRHYwIh38c884li58DN8LsecQYfg6dDrLXhnq2DEV
exD7mO32PLKDuEN8Bsb4uVAgs+gb79s1YGrxd5OoQucmo97uJHZnHX7OzJFEBPgrx6V3yfvAjlxD
Uxmi03H/eqORJYhuQC79IhRj9vOl1u97X3syf7JEoweFYkySF7vkh0A/gHLKORYTRp4Utl8+GRUS
8ySZUgV5VEhITNRhau987kyLcvOrtYWJUO4h+56XXVf/xKX7H1PHqp4CNxjHN07TM+ARJfmy3Cz6
VKxwf4KEE760Pcu7kiiaDF22pCqilNaHDfSRNxSUQSjQhFD4dSfNrThn8Nx6EQljChBxfXQjbwjN
e/a82QvqrTiv9F0hJUG+s6seCOxtHcGPqbzp/MvT+JgpQDvxXaAf3cVxaky58b79Dh6cYRXt1cpH
lrDqafxnNySGZMKvfeEnRJ4rQvA0UkPA6AYNOUnJErHq9heUXocBz067FUR8RfFA7PCPpMb6ec+m
axU7OYtoUSfP1Blz++N3YHygFgaaysLoFAkr5Mc4B5LmxN/qSN2ONX8xHvr/CDP0m2y2p0IRpxzw
vbXCIaWzTOyGBYmhtsOhlbVyWkWtC/3a1dCC3Glk+Fz6vYAqcoGx9F3K13oUbEk+7/gF1LrrWTLl
mVek3n2Sn2yOODt1GOONzuJHxEIM/IEGFbL5bSd5yVkPBKw0GZa5QWQM/JRMELbCsJ4Zc6+ju/ur
BlzHor3uFnd45Go9d9P67FfVOlv53ShKzVuSfZZvId6kY6eWcxnqJ3ktfoknSf9SRt76jgZR8KLy
Rv05QiP4pU+GWXyR7JvaaHzSvBhax6z9YGIrpEPWKyDP8zJPGblqmj2q/4x3WpSGVt+YCUC/pg1z
DO5tIoKnXq55B5TCoczWkBjQjUsiMV0M03LI5vzP9H3/Zle8jMpzceHKTSnbqIaUc+ciRVKaOgBC
nkphVfzVcZQRgxl0/6xiwT+1BmoQJDiShEH0+OEi8jzgyTEhBr/Se4k8TzRD154XEC6m5UOEw1GL
+uQ7PIfCFxC0K0oUnXyWHYWexFR8JCY+hbUPiUmeT+BzZyijVYhSmEn6rW9D4sjiXK477YzJnf2T
xnlvtOOLM6HrO1bQCvNaz6slbhU96mNQQHLWs+8P6U7rM9VB7QdCdgjbmt1HnlwqqzYL/YvdTAf/
PrHMmquLPyAUfRmWVKUGdY6K+KSOsXeEBlMtpWeh3O7XbbAOdyhY/23GV87Ggs3uE5bqFKNWzANx
rQ7iq+EmupeNpOuBhUMFRNfjUuQMsBmcSXz0Ure2c/2fQALgnFaXVYeGsDG0DjyzIRYHIxkKL+22
N5+qR8aR7zat9drjb6qrJaDTHX9gtkq3OpD3yK7dSr0oKex/uVOsEqbQ/ldIeL301FxDN33/VWX5
zqNYMnVDqtrRgip+gi1ewOOXzyo/C0VAGdjzc0rlo3WxqKFPhHY7/Dfzk/AIdI1rjjhvKbHaJVD4
hOHTlN7eSZ8QmhZqtuqqWmO3u5xWfsKrh6pxAsJMsYeQvKl/N+PMKint6rmzezg7s+2BSO7+yrZr
V25lfgtWHCrkDu6f1A83VCepbg8IhixddX+ZaTK7it5BhvPjYif495AkOF1IUdJMhq0UVyS2Z/s/
Mnl7Emj/zflOxMVMov8CAvxol4ta+d60xE4CZiQbAvspfVvN56vaQlxbf1KzwgHgNYflfhuDsUSO
KztlRDqBxZUbUScx//dIaWfK8fITUpCPc0i8rfFj0Nubc30Cp/pdq/tGuezNHV5hZkHroU6/NlZH
r4YpU+DTyT0gdOLaV+fw+6M/FltW8nOBQwXMieAxhArZdnaor1yr/99d4Q2mTSVaYGEr0tbK5q9O
CmXaUdeTqqEMIKTc9tIQg1Q16b5r6pgyF4lqzOSl4a/HifLd3zNSkge0/64hC6nYWJWIUx40W52U
J3B94uugSqZkiLxFs1Pm2RwQCf+tNp2uMU39s5Sm8F9mdOpEMPoIU/dlwVSEvlrtvg0bJc4O0240
KC/IOSG1890/Z4JscC34z2kfE9u2JZoe0WEMYKOzkeo3zh1tguW7XTiSNukRibwVtV8Ymnfwjf3B
lhylthTQNqVKrozusUegy8WKLmsKFvXAf4rmxyXQ3C6LntX2onU3bjIwv2ryFjd7tuniAxaDKuKT
2daM+XLqujicuadOojL0OD9aaxySim+1j7FBAqtXwkVEfMAXiAyoK/BuzNklxWw7K4mpmNNAADAU
QMiGib7p36icqk6GRFCLRQ354gXA6wDovT4nkosd3N1MwQWiEvJB9uuyskxut3NX6LfjAnxtWgpM
8diAPUXPwcMJ1mmMcB0A6GZQSwAn9kuEF7H62EjntA/cqMtHTw7CWyWgynfyCqcjIIiwOFR9dp2s
CflRv1+HYGX2xenOjVemz1Uj+HgPbigkb/SkCe4CjN9oLikWr26k1JBc5yFBiQUUIIfpMWEH71/E
UDorFBxYJDalKGD6n1lJsY62EuIIb1xpdElugf/vIB8W0Oy3cUwr7Faykn6BuNjQelqDfcUVMgMI
w/qhnefLlQGMYIXj1ARr3N1LlZ2yBP85GatQ0jyStB94NNJv5oxZ8xang4bplAnJdgSXQMoiDeO9
AHnkhx4FGs7bgdVZU6LNpBhKU5Yvf2joJZm+iFBwYeX0HWB5+mckVytfwYS32h3Oy76jETZ/RofT
u4NwTaMgN5OoTNlX6cadVxyecsoNpGeTK15mrtwm5V3g3SFB8IAReXha9kLweogdAos/1sNvYzG0
Pt7DS45qii8g49YNEx2P5R7G6fA/72A/di3xrDktTlz6d7CPuheUSQnpQEx5OFMTG+KfmqfFYXl7
3MGy05+DcuKUavkn7L786s6rLD7MX19le5h1Y6dRb9CvX5fboeorVxzuSpDsvNxpIX5gPFdfw1C0
XLqWa8JkbfbD77haZL9OHQB/FKIMF0yNeFxVReOjvY1/vgZvIhHkr3gaDXoEvo18uiyMETBECJfX
wjDqlan8g8PQLtctq7O/GgfKgytG3TLEzsMljeL7+FXqLQd2iyPguklnGAQdPKtLTel/gWXitpwA
r04VgN7dOfvpvRzwwQrvyGAvd6CaMNq43mjhiI5NjeRloM7MTqu/+aIcB07UGMo1LcBeCxiMmiA5
jpesZAWra1MxwnCOOQWzEIysM7iwIA1751tLz4ztgeKF3gBmi+Yx3RhMUpnLg2qBRGeL9ec9LFeM
0JHJKFdJ5PkTtx1cZZ+sSq/CyV5Xvj7E5j7QbE5c6FkPPgfE6Yn4s+pgMkshzu5+y+y3bLAo5p1S
dwS6ZhQVAiB3xKXHJoA0wd0+wPe1GdVCvRzBWvsf6i7eB1WS00kHaV06dUJUB2i8hirzQGA7SQLV
LspH+Vzd1Zole1vbpa7U4iTDROOZV8p9jhkMDBoD01kTlFxda+nGcyuh0OApfE+w0XZlOpXDdSp7
VJxWH0GUf0AM0G2ZY+E7KorRAvIR8Vbj0SnMTZk70dFqaVSOb07CHmtxxIHfIFu1qTVSYg4vxBg/
wf1iJdAg3KOTnHMo4C5njZZu/sQgLmx1qWpkub+pnIlbnTXzvWeuIGRD74pYvEyUT/iWlKHYVvoA
JNQNz8F19zfkEkksqs1a4BKQSu4d8uX9uTr9Paz16cWHvq5GU2X8kMF+dpAxoLEK+RG53CwLsnoR
vSeuCP2I0B7uXQ1u42zCEX1PdEYpvGoEWJRJvmFssMSmWg0INX20DyrKkY1fODvLLEW8DFkkrReW
kT7SiwBT75cqBVoe7WvHquNUK4MupuQBIU4YWMQlrK4r/8ima8lsiR4kDEkk55YHiCyPKhT3RcMB
COWK6l8YBylxqJ6N5dGl8SFL9bBNMD8qPFDM2JR0x4t7dnJNSVpvMM+One3hWJfmVydl6kvO4fFF
Or5pNJEUNHq/HEPpK3l28bGqIQGCuYWcwtv22gObsnUYnRQyQyLTtriUfeax9Mp8kEFiS+WeJeGP
xsWve0wGKGm7LBjN3ytLuhrDLw+NaenRMSuZOE9G96tU4MKfeshgr9/NbeaCZxTjRWPu95JdxP9r
19JxcEKwWuWxGsw3NL988DP5eR+M/B3dV13GydkAz8DIzT2PNesNDNc9IlVsb3zOBVnV3oL3IfZs
b2w7YwAupzc4dn8nhuQkGfteAn6claxBaYnnGzqKQZ8H0h2EQ9QBAoWAiHsADUQ8ldWr+gbUr2lM
Kh12MzvbWG7pLBQWn1/MaLmWf5N+aXm72y9Zn+2EPrbDUnLzyK45RXxIJAJ/uiD2UvrJS7uaQryK
6Y00wCVrn5nREZpgx44esG6wEb05glc9TFuCNF2NL+8C7I0xpBS20PVAiZPAtwgfy5p4l8y/ea0R
4maZACugKH3q4293+HugcBjDJ1dWIRX7fGlg0pl/VD1bqCr/vwm38ViUz6Fo8M1CPQ6nKHZi4CQg
jlZKJIs89lNz16//32IOBjT9RNZBoU24aM618zcUv9Ca5ZpbVYct368ziUz4yYHj1iGsZLatInWn
10XYwmzJpCyO8Tj4S/pdQUREi3RLbBgzC0yl2xKUn+DGPPc0iUlydzynRKgoVanxwyOP/XOkb+/S
VeJLzsXwpXRwV4ZEzwTjuJVh/qsEqjFXYXiZFoBNjQa4qzfbs09doGIscmdxGlkybBgRnZDGqQeO
Mk5vC6PgjQ5TGN0q1rM3ap0Uo3KejLrsAlSzc5y8z4npPLqvYH8URLOXHwyUXNEV2yexfZzaHzIP
U7ddB30QQTCatCAoYONlXL61Pk4R8TIjcSzG+tUve/rTq1rWrUt7vsIAHId47hOs4dgTVY7AG7lE
/IuxI6OJwCDA6Ui3iPz+NV4LOzhCjbj4SBgK2c3n8cGXTVOI5YSOeBjr4jOzAuAZZIbrwwzSUQLS
gv1EcUIO1MYP2NwC4COk1bwu2PUBMVt9RuRr70U35UjRP+2gsOaTJoSBMoBnc+TqRj9zhb4b1Wls
44kVtsi6QnhwWic8hQuhA3SqmGtpXE31ZpRFZdnXnG5Fe5pgY8Yy3nxh+1ktdHU45vKD+4gKhK09
E/QmEJiWShkGVQVxfkfUFzlXkTM70xldi8V1KRhB2lyjxLv4h0OpTddNNAsWb6stgUHlUBUqzDI+
uESoo8kGHVQYegyCSPJiOwyvi2ubDFVQKXqBylwbLmbZ1UFLWUC1o4L3MORWmOv/nBsv253vMzlH
+xbXYQ3I4Y+osFfGKwnwa0HN+Yr0JXBi0XCSr7xUOtbwIkCZUpShjCmMQ09UEBIc1/9HERyQvRE0
B2sfcS6GPCYnHhlWZIUxLHxFJTIB2fQMOuMJKyTu1mMeQIVaj0AvaAmV34Qx4gqc8Idda8UdaF50
kn4Puej/QkLdPEcUf5ockg10SFfVTZ8VAMNCrwMKnQSK7qqCIuF5Y6YyFjWjA6qj6+RHbcZ6Bz7d
574Xlszfs/qJw/THmWQLTJpNej3LbshaMBmKWYuQlNnn3ZXeOJBkC0M225hntYsPhatRMNilDlvw
Erl24HYOhtYC4xuQwoAVuc+EOTAoLjH4pGBuHPTwOBN1KclZnF0ArtEpJJYKRTWD/EyGB4xAiuFG
o10NaCqwYOo1YjB6wvmFEkDdBk0Yvu8MK+kvJJNDF8VGJIPsr28Wj7J1GPxP9oHPJ/r/e9hxwF0v
kEVhkD6Oz6K51YJKahVGBet2ZU926B5PP5TD01ukfJH+yAD+dT9HOWw+pwE7JuerGc/tzpSFc5H4
v1xd9uOUtvBgY4VIKJ7K9xYKJuIxoLsmDzW0GqWenzFZRZjsAOqUIyb2ZnrhICRZvGD4fjM9hyiA
pxkHU9eW8U5nIuSHl6+sm2KTU3+MyB6A2GgF4j/O4Hg6EesV/CVmZSaoxg2hKRCiC6LiTDcHjEio
g7VoI3nRyiiIwyCuFioWKzzXoqXl338vh86mH1e6IVxO4AuQisFbJCOJJgBVFfDP8oP+byuH/eLR
gAkpmvC8Hk7SzAje1aUwlPB+tTtZqin4U0g+lzT9rg3ZQH+RjUUIgt5eaonKyjdGNsLX3D9n2bkX
yjnBiZpLky+QFeQ1qZ4vSV7MfN45N1CF9jfYqMPQcZ2g+w8qMjeKhlBAqCasrVttOhfGlDScuPUh
3Uk+QJONnOfJLYblJ7lymr/DOb5R25QGIobOFE7y7FIzxMgIgDUEFfAvUWtXAUwoQlFCIU10uCUA
emYN/Ol0EhUCDprakpuJHi1B+Y/ukGPjFti1WDMQXVJAy3LCYvTiOdFPFsVyEnboUhDXAt/bkdqX
rnihBezsXwcLE9ebm/q2Y97gbkzUsE+JJu5+eXh8Ee7SJ4lo9+ph52xxzP0gMSNDnYJRO9/4J1ff
IX63t3iONkwSJEDfVEkwQmrZfAK30Hk7R60CO0pTycgnODz2T0okiljG4GqFWKBe7sMOcR2SzUU1
fzjKCMxJxwQFblu5RZHxLtPtolTwvK1XBa9GKdoBzJeBomaM0eWJE80UjUIcJD6XuPEpDPHYd6Xn
9sZCCTWa0XNYzB2hRNcxlcgSBKmNvVzOigNS2h1CZpeVRfDDteA7Re5yDesuBmPl/8Hf9uTqyeSW
50R8Y6mJ61yOptOLHvGEoSIA7zvkxIs6IK3NBY4mXyLfFdcDaKXABOw1KCxZXWw+96E0WZ/nksxW
tevNBYxyXFuOHQvSLYrcldGlQh3Dm+/tTzl3XREboZyNQRV/M1Tyc38ok2jMGdJz+WdQoGiadSeA
nV55r0PU65f8pUfx57U5zP1psJ+elim5FueC6Wly4rnLs63+DVmPkbnsUA9JeTTjkHi4kKYpE9JS
04QoNKBwY5yLfDXhes2FQfkU/Re0nfiBM7STLsk2SVFboTf1DSmOX4sTFOwcqhejUvO6TdXqf4RC
tnZsEZ5fl+CU4UgxtE8ncKuqUzU9Fh2M8f/41hEUOV9KBDYOxA5PqGB3hVfBR2BVlL1mKnMDzyKM
WQoG89ZWtZuMc3UJgO4nmruy5ZKZz0ERmhKJhxefttLkVfZG6wbEcQguVTpQWBHw5C/ovgAoNjRO
amEHjEzzuZjwW1Xedu0PFFDj9jQ5vS1py9upQFprRhzR5Ca3g6xPMn4FLRRlK8S9ZS4/DNT1ZP6l
G9umna73Z6lC+WPS+7N2BQ8SWRlDunaYRadG9WN+R2l3kEwZ2GGVxzgKgsXm4AtxX09xIcDoBVmY
15TZGnyRxH1P3TMV/+OqJfTD+cg021pO6DbpnJhFYkivc40bvMCJdNHI8nK9ysb7q0PS1JkX9N4w
HkXtNPOy2M+wDM0++bV9lQHNrrp5vbupe78fBIOvMPKXOHGheGCgWjNCQXY4sbxJPXpmrIZOpR/x
YkvWrDydrepyqDUYRn9QVW42LBa6kaCsqJpU8pwl9Rbylkaqe5pkTi6DVc1uPW7Tav5sVmqhXNm8
RHd5ow0m67LgZI4AeJpxbenFRdnLZn1rYyxZzePnFTzZPcQS2pecHGvkJMeoFkM0x5I9m+Yu1RgH
trft0ut2aZe9p9CGuMGrqyFi9xabfThuX/1rZI3xN68YrAgdUikPdMmgVJ93J6YdXBobjE/p68aR
NSTWxtjo+xgrsox4kXKcZTNs45SB+4/8FkWtJsF4sqLwBH3wrQ37gW4qgq6ihsSSUiinvZL47DC6
F6TMS8cYXr7e+fs/TzpIZMBzTpTVJglrnw0g5HDsznkqLNhAIogBTq0FUTVA8HzdJ828kiD51f+2
KBYIPzjGQiv+UFA1CgTQdHEasTAmS9yHVaeHdrhsg0EvxPWWkybPJ6obcwFbeknpDuLLQabXsbpO
2+kFBKswtnzHhtERG9YigVhJ3lGYO8l46Ks0nHnhesKasEhJ+nxU88x3dhBCC++/h3huuUl6qaaY
hY3FVzc88MQ4FwK3PJ3W1EUhOGdZpr5J0kqswzJxOWpYi2hX9reX4n1e3m7oym+gRG1YPSwIDfTr
/2RYnMqhKKXL1WI3skWKu7ZFiWnnQl3P85TLPMruXTjemp8e7PZ+Kwk7PjF5o6jZiyQYN0sMn1sw
37gAp70XrhqlyHVm7Uheul8Sf69Vqj+Me9+Xb6PTvRp27qI9eG9Bra18ePaVXJgJ+67qpzpGjFW1
7IQrwicWNtPeXXyf9N+Cfsh9MRVAqDwfKxDKwWC07cErSscJw+9jRs6tTJjA0FUQ+ZhHjuxEixVW
9PEY1VM8ACqvr3M0G3+LfRko7y8rO3FV2RfKg2uZi5oat5r8swaSEZLBKGrgzpUQudK/N9WC92um
ff8h8iYKauZF5Ff82ugmhyZ7ARXqcYPcmSHQWvbadXvp3ErqEbBbGaucSiNz1QNcDcNhc3ZkkvjJ
sK4EiykpxkSGVj7qpPtDZD39UnAca1wegOBNAsgjZXcRb8VdpLugB6XcDx42kI0TmplGssyUqYft
tpLxaEtRRBdTUkEV50fYJOPNOJHut3VGW090Nn7S4Sxj6FC/eAIKZT4TLbhqsLIZ+hvRawYxtzA+
skxn1sPGJHQMxiD/lZaWJFufmm90IsW+V4IBBKOYmEiTy/KDqtAEFRU8lXWtzheaXtyU1D7Kup7M
lI3c6SKFjUsoXGpInwuHe56r9z103AGIS2wk87YEtUHpDyi3YakZQG/Vy8aDVM2UP19zoN34fdhc
GTXIogvwqKAFz75STyALuY1NT/mEQSkootXdfrkviRdyfz93z5XqRgRpuh8JiyBqLk0mvd0tFS+m
sRjeAdjrruq87gOcWS7cFJUhArf5D1OpCiqbMaxXyyttHTNJaO1M9v2hCJKhAuIz9YKDxyQOq6so
NkUCHqpOd+qecsN9eDEsHWHOmKX7B6dstTffNNKLQYJpoJO+Mn8KdpLB1J0WsQcY7iW1LqC/lT07
Ww0r+JCZGsgPpnjgxwxSanUD+xv0/Xc+I2rNXEa9hbv6CrdrnLKphMv0xJ5v3hxkaIzB6qcr+rno
gXE7oNMMFysNjDr4IMjQXLCm8ntB7ZBv9SjmGwz+o7Z/8vpDdodyLLbWluL2UfDEcQTkEAZDRFDY
1rXsrH5VLoa6ljGY314kJ+qFmK2BXIoUQvOG/dXTEXpgX2XebPZltBVjOOZZGfynRK7foBqbvgrR
f14jvz9mdvTx33XSnVzGgwN05PgCecRyhhKFlmrbjsv2lKTp2sJwBbN0AR84B5HZZY7kp4/l2h4S
v41bftpKL1Sbu5Cl9ysi3wZRaAcF7M/sJA2asyy4p4bZA6wbDpm3Dq5oKhXiaFSkCLx6+AcE07dT
Oguj/ELYgzCNqLY92IrXf42io7/SZ9kXSxrVPFlA0S4gzvJmNafA9KE1B2FeLP+NkhFOouzZzqMU
jNpNbR+0F/eRASP3+t+TsqsHF1zNAYsn89qmZ9yJ0dsQlG6vtYvpm51psWhG8Iti01jgyCAMafgK
7nQPeBAqw1iK2uyOOBoiK384DZGT95OSvKHG8SQ3kKBHJgdOo4SY4Tnz8bMeqM8lW2uPLt1yM+nn
MSkCeEX8ZzJ1ln4sH1NFDpjPh247VPKOYi+4CCGh1DoEuCwgKk9sgE41i5NvAOxxiiD5js4B2btq
oZl3cTPHuDyUSvFIPn6CrSq376vtYTV7eaZxcNgcmcSNZQkIA943gTg8z2BfwKMOHBsC/bDs+k71
itQckrMr2ATTCuHaY/cKzRFix+8MTVEU7Qj2gvn+bHWECZ/W32BSLu8MVAE2+8lVGTD0UJr2Tlzh
GVY4NloQ2Occ+C9abFF4y4iER83R1XtejIyyHjj6wuJV46v6ezvQ33Ov5IERmqWhXmCgCLMMcvnw
EORATRrsonLD/iWZSIE2yQwKPOVhYB9mGUUsSr2v09DGfPQRvRBPU724SJ1e0me2R1Axq2tPLZII
KIsOHeA/GnDI+IesuhnwJ2mFfDM93l5sMWIxtSYG3Km9k0IdKSeg8SjjYTqdkfB4dbpgPvd5UX92
lieewEn8LRLs0XwJJcU5/3wK355gZ+Kj27bNUhsf4j8MvBdqlyNBgeFU96cRojcOjaT6vSwBG1Dq
cR2iih1cdCY9pjfsoCVA9Em1WS+DeTObYJMwwh4J5y6FrJ7VBLE0ghQ2E19orXKTSrGCEGTLB4EN
2xVzRXoLfmYFMEPjj00teiqmw9l7lzhL3mzTtnDx86Dy4MPhrHs8Ka9eDjayPyykFItQumzLn1aE
LtLwfnYO/4zPylcuJAVvx3L4jyFda5WpPQ39Db7cLY8b8JxHj7XKYslYAyguvQDKF8Sjm/y/fZlQ
iwrefkHKOikC7AuEnvwvg4k9Q1Nki95chTLH6GyRXQ1hBk4YfE2XTw9SlRdJv1y05Wkgv4mZNnda
IK0PwT4i7qqSEDWvqyPpbhLM9IrB+goRwZwVudd6g2JaWSyc7PqcWTwgJz2DRBeEwOF/N9UGOpt7
0N4gyIaVTExqjUZeTei7nPMQKvDk4yAWhLrz5Ym2ymzFw2b4zbiiAPxnf2DXUQjHrGCju0XpsKnA
4SxYF6JY+f9JhVZJ8otlNIZGFky0oW2vC+rZ6jGby8/DzX5dLxgHM8ztLIRm4q7v1S2hezmepIAQ
ebsFbZSts7RHUk7XvTpmuguo3dOyTXb4Xlg+wq28jas/HsuDh7ikYdIj1Lv1cqcA8j8C3JvpGYM8
MebU2gQdsMZbycEp2Djs2tGkDl7veQGwHFK4FvtWmsOMxVceo9uOwLiod4aegwrusv3L8jt7c47y
W8kIOg5XPwWN2+O5QC1Nw2+EDlff0oaXHBULbroDfhKXZey9lBOTGg0jPPS6lEpLDjD3i4nBpGCK
iFvWvsDFvyDz/DIpPWWBBZIfhzrmpPIcCtP0cauNgghO+LMTZ95Nge8chKCqnsiOR6r4kV4sJBxH
CVkGkvBAFicKfwi0r0if886Uri4bbiVfSdeNAJBX+fePav1DoshO4GFT6/c5qQ58KihVTTdP+moj
2PJifpoU1KcJzSlJNSV9T+XwildqHKn50JMs3CG2CsGxtfrzPyVE/xpQnlgJp8A0TD+xyrBgGhqg
zpMksvT40GgkdJw+/WiVvyF5clR1Y2Xig8AaqYq+KPabdux3cXM2+zKvY/fMrthh6iq1STdpz487
a3lQgHtXFF/9r7mIUOUBzQvJlATkOo10k+5J+2/udAb+E6f6jYyYqZkRXQQxPCnv+XJfY/xe60TW
DGAzPEFABMWyZE7ltVlFzwLVERwD1YoHirT9acivt32y5jOUg2FCedZgEtFyZmlqQNKE2ESUvYNA
n3E9PEF3/NidOG344INw9P6lk7cMoAbD8V4KBtjyfGyeOZqaLF6rlYLF8K9ppE5Vh0gbzsI9GgyT
bbwVzGC2eALLIZiv+ta87Hrxod/gdsD8Ksu5pB7DwtB7gkDbTGbm6PFSOjY5UosE4lSWlB8AJype
XK7mdEMV46Xxb4m3dFhAAmsYscyZrF67EmxE/FNSMMUYse2tBF80LgYR/NiG+EhMIXL+rPNXf4rZ
dZrwIdXiLtdyMMKHbz/AUZN07HUU9KEWOpSzTGUShbDpln75w3KANPfOMBh7OdU9MhionVeEZxOZ
6MsP7KZnOPKy6YWRXfA/O3+KbrX/wx7RDSnFgvGr1od+e5uRBicvDaaAJDaN7EBOT1bgmaZSY1kP
2EOKPy3F8Tr3c3sZjTtSEpaoe/XI5sz1YZXlBlu81L247AcQAtLcZjZN67jDUvs4y+q1TY5DTLC3
foFD6LtE7nzoRxvRc9FOs+JnFIp7/+alaYM1blcG+TstNHYtiVZs0Hv7xHt3e1U81U4seM8mYGGo
wu9nlBgQgr/YZBfAFSqvgUHlBgyUAHBryUnatzJkIdcwy5CPErZ3dzxKJWmPwoOwg1lge0hZOKuN
aYuusIK2ZfMgNcm6plbCadQ8EsalCRdXvbL0ceIMTi3jqJVK3qcplu++f80nzCFVGe5EUCdBHgf6
B6HwNxkEwRtReKuBRVmraUDVErmndv4bJMwMUbu3URPia6MXhGDVrECCIbx7lp8UYEEICMZfYvaj
MVTAz7fdSpnc4qvZRISBfDnFklK9fhYY7Sx7gsUPBps+fpwckJHotqQ75rsgdyY8C14tkZI64wgj
NrIXXU295S6dzyKJ+T3NBmO7VG+YHuTkcanotHK79qlTzvipWpdydQIK2eY1BJbeYucorvWQb7sP
mysVJCjlzfiuR2X3nBn0J7XnYnsFM3Oy8qlDoONeWjOGGuqQaZ/CgXJNGg3eVNqm1/y40ItxBWLF
nBx4AKYvLNzzjyMxFlHo9VmVs4phAzuFmLvs5SjSdy9Xd/w2k6GdFcHL/D36ZZW+0E/JE5YgQrai
pmx7Y3vYFstaG5P0t87qPFxojMKpZwWyhD+E+LMWJdTIo6KW5j4VzpITw/S9u+ZwqmSRD5kzVLH5
YThBUy38ZAEhef0bBlDnHC+MT90ijSHvrPmXhPkD0KtieAKuBWDN6JpKp62z5tNZFXvZ568ftEZL
ADQvAiro5/sFL8/ZORZJK59fbLDqAH5/u8j7VA2J1anoc+zC6LgT1aQ4craS6LT+LY2bGxskH/ST
dRs9RIhacr2cUYF2IgYRJuN4DC/jZrscIn8l20xjTlvMIQNTzSuXsugETW2XOSVkHpCb1UNwRjTq
/AKIOcSqDhC/SZbmg5HWrYUr/5AZTYG42lPgDp0+wzPe3Aakz5XgXXaS9A9Joh09eR7wGe25Ks/i
T/ALex1JGM4I+PPd1z6ACngifmOQJeWEZAcr4vLqe69HzpirvFffTvOEyIZ9fo2sU5cKrcSO/drw
iQociJV98LseOmh2mIjUEWikC6iHBu7fAjy35Znu+VjHxShjQRG5uDhVbglb/Kl/noOMuhJXDu2A
uHoUeBUg9EoXar3bCfeUIg3AuUUxGWfEo7m6Igr06WUc253snPkQ/gLHbNQlsJFCsXWcGBzfBqmh
GAqB2hljK89lgjmDVL9j5WcBkAjHD+BLLp32qvzvFZ1nivyS27H49Pr0o9uf3TTGDYleOLjH0zjY
a5U5zRrTgegMasDF4qJtiPONVUFOVACveLtx2HrN57zPlwIABDoOCBSEE4LpKbJ36eiwE6XSGTqa
a5SLPCldttgYdlN0JoxAQ4TBzFApjqrrtLQ70TAKrGzwr1GXxFcSDEoIglyP8uIwk8JjqnCjjsMr
CZ3ha+59qRZHPDeMOy7zGXvMaJv4aZOdTVYV7CXOjk6qhHa5iovKT272rTHbS+jHh4itRS7CHIy2
lhg2VciWE+iQH4RBlh3m9kxKSz+XOtDr1Rx829uBONfE97NdCmVA0T9qOygFwJ1s5x0auHlq2VEX
LvmS4Yu5bIZ3ZuXRCjSlDGMNAgWa0K2c9kc5g0eGoDlR0Rr/0CoQdLwKkkqypbq93xgftb1ZiAnH
QMI2py8bRsRPQQSMqMaggmmcN2Fo6bhcWT4/qV+z70vYqEt91uu5K0n2foNC31R7cPq/f7JMHWZl
ianPB+XVECTofPwWp4wAHQ5ruwOIke3Af3TNfhSW8HEUKdFtrrN9tGq8BPn/pI3DPLIOUXdK3edu
QkryDXHfLRdTLsmY1csVQ1/nEfRG96ENMafwGJqWLgz41Do4XoX4NXhkkJEi/T1dw+shqmMq7lcQ
31q9UNaG+HV2a9ICmywmK4mp7fXkCBS4auVVy3hbkGh7OUe1RdB6M9gAx1KZKoOxMK2vl3FgV1w6
Edr6kTQHAI4RzK1TM94FHUDEMGNli+1HtXpWKuxmieoe/nwYlwASmDHgYwyiot93p2IT4ATHgJDk
xbPoMzSWtCw287JIjTCzTu8Q/erElHnBuzW11kHI95LKHXf5C/0J7F6AcPsailOTlvNoB7upL/Jz
u0gfewV4EMZnUIEFcPRrKmbjP0hOI+q1COIEEgsrKckXas4LERUQ0U3XlQfwrVIVzds+p/K/7dtD
BGeeVGUnt6OUU/u8Vqu4W5Ihs+Gae0BOG39ZTnWSh7AORPpP3pgQaPlW6Xsl7dO86l+rO2Lr0PMx
Cml2Q0pZIZDrbGpUHzbkf4EcU1OoDvxPzym+xXH9gl9rccrLHpZsr5bqKmu/hLE3+UrSOpeU0jod
6QuC3gKPEoYT1T8kZAGNyig9QsQdriqEPWa3rMFZg+iDAbC77/q3K5QGyc/yNsPpWjAoc0aDNYLg
Bk+cUSyKhjU5X06QIKNWBD49Nc7fTx9pgp6FQ3JMnPikxrRdwwBV7t2vJoZTFWEcCI1n+C/XdWQF
dmmpYw9mrtOvM9J+XtFr/ZJM9PpW4MhzfzkDs5k1+woOY/IlYPdElKeSy8IhhMx8yfTBIa6ufAbF
kGD986uFAs1kimozh8GPy/WN3ZT5FJ+bRb+G3YA1O43joEp0b6Zu+zzJRlERN9fXm+OZlgolWVyA
irfL6+EYR0tJyAFPFblNiMFQUJRekUb2GqQ5Mi7wSZ57rls/B45nVFKAEufwqZjp33vVMJz+buFz
VK6I0A141lOJm5TtzKLcE0YxtvO9M9uYFkzhTp8vJEjjHwlDCK6fQxiSbnlTT0ibfO1PwSWKF3tu
F6gJkAdjbPshpqkaMxiF//v3/4Cy2ffG6PGwrq4dyzpXy5dMNpYMx8//CtYG9OW85cK5ybEW0qH1
MFo3p6forzgunn56YfyvGf3Jg0rc9JdHp2OFs3Y8cHzpyebnC6Sp+ZIg72OxOzEosjmPeufJUcNB
vi6LIyL6HAVM79wWhQopKDao9N6G+oTyVUJFbz6uRlPgzonxP2vxJSMuAvYnfUbSxzqwM01mh4mm
k66jl5fCo20U+IiYNsqAc8dsLwGoCh/oY8Ej2aZ02yCLdWMc3zLrL0r1/hy3+EiiKb5UohYxpWqO
Z2seC72nxbTLLIgF8jsv4DKoGEljR46Yh+Nc9rWaVPsKTdcW9JjnYdIa6uVfIPk5yCyoEe6vAxZU
I3qAY7HmhtVomof5kP6Ky5W+/8GExM1InolbQqTRlQLm0cQ+l832vlvTJVCnxACl0cxjVNCWY/Ra
cz10DJGovdHB1SjqYBbw+adZYE3x6EU2aGFMz5FlNyrSjwgmB8Tyncu6KIwvx5ecbaEpajcrC7Ce
cZ2m/MQaaBu8H6GVP/61zx/Oi28y4dIKBAEVHzLfGVCGj06evXvYC2VASOMV4IgFy2sd1hYJLZSd
8qv9Z+0f2K7tlwy1wNY8G1ifZTVYV3YF38ZS4JEVMmZUo+3NylrJWpdbtuQpBMSdbrO8u+zX4Twl
XWJPiJE1XGNcestpNQNWOuJe+zY0DlIG2tLB7C+oOaFRJ2tDMgPY9JDI04nxSfS4SpJDavl76ACR
nAL8J2yodOyu7Z+q8CkH8XByE9ZiTi1ugZoCITvnckJEWhnUUVKoEWfaKEtlojmB4qQ2Mu0aWwHg
vR2zZUG0/xLNS13BFgEnGl2kmP2porweHg8QhVGvgukjfNsEqW8MH+qpbIAU8HfqGSC2ODdWjbJF
4VVkycMEadTQYg69hTRX39FKy8y7m1OFywUJIX6BBh1cDcw5ju/gtiM4Gj9G4WWhqKSZzyy24nOp
VIUy4ZHUuXqERJOLpKfb8ny1Ag/jDPrLYC2FtGF6CeIc8NBEYBzB2OueyYIgGywU64FcmN8k1yGo
2CPy0lrO3tmewD8yie373BDETyxYA2/KncXkLo0fGx9FHwOaqxmWccOlIcnY3WSUf87VhPHvfvbI
Mo0yQs7cU2DwhlnxnTTEZ2wYRPemMglKW7wsu9ZRnGK/LydLewOTf/9Vve/pRzCYbFMLtA8u2obr
eb2mUz8yiwVQUbX9URw7IjSxS4lQc553jNVn0rodsBgRTqhgKnlLFf6+y4nfEqHnGaOzTCZlr0Uv
jMEqiagDsRMQ1cysuPGkWxR+iRzI6fdqyj6yn2NyuGhq2/FJV0U6/6U+LfMI1h5NExG6FfuqFjBJ
9YPgAS16oitYtKad8UPFQs9k+5+NrOLrJz0uhlSbhpFNpxj66TwzUNT3uOtQqKXsvzYjEThRZZfQ
YQ46UvoyoBMuiIjZNli5HIzJ1TZzGoFxQ9/MTmhyVA494Fmw0KWnfYDMIcjMLgQkKIMsBCCI76sZ
M9ZCH9DHa86S7qRaqEeIdBR+LanalLY90JuDv3NWZ+OKfNVtz6E84WE8GaLt+LXJNpyG0UPp66JP
yjiuQbhD/RBhK2sWjAmCsyEQb6hn/DNL+PC8CPBzLcPgMrX7pc8hWYGSrbrGr46h8bnhsfSjcQVF
XdkJmkjaLy65Z8TMBpuK4LySRR88LFThBYI1aWZ2985AFNeMygIlR9RNMvl5xPqLzBpC1naSV/vY
VEcS48EKGC2GkOGvrfE3eTqqs8oxGkQlRrn+mlzpNaO4lnAzTsabZV89dUESBu60f9c+Tq63wUlo
5G5+XNawK3bCGNFAAGGMuRIDoH620y2yyA4HljVQDf61gywcunQzWXssgIDNZnfuPix87j2+iTH9
X75atH9cHCm754IjXeSJdbcsy2If/H44Pmt+eEzaF7rs3FNZSr4Y2P/esNWEriGrr6EEcw+Tu46n
qQVRgzUHq1Ad6XqMG1RNhUuxtGTE29hW9C7wLR/IKtMrzJjeSD66WGv4L+vqtQoGTNMHFPA/ovPT
9YE4p2i/Tv/aJ2DzXGWuFQEeQSBhUGfbOBkxfqQeIEAVXbdzbmPPVjlUvWdeLxSamEjxE/b+3OpY
5jr1e9FtUuBnhoXv/MTvF4usZvCrkzF6GACfto+upjRrStKJs3ns4DmuD8+umB9lcUHi6LvoKvZH
uUAxVHfX7R3c/vU7JFEKvbV1uAOygslHLAb5siIvEKpG5j0cLt8OCYQ0crX6hRMburVwW0U0gWNr
Vbk70GJGVKpNcFWbnVm9PplxXxxtlccByTL2Cfw+dCNrEUe+urpiCI/KRdoIT+XTC9EJppNvkvI4
NhmjpfNJmOqvbYX61wwxJudAd4wiioS93UIQ9C6kFJVL/xoLGzzRsOkDdeJdzeTinXcIu96gPpYe
cHvWWsN/2jE3Lui0qSXBlPvvcLo3dpf4qYSuXvfVlsascYsN5ZUv2oirpmtpW7+yKg9DM26+0Dwp
p7tEodg7NK5J9SQR5OSXNq48rqGqjZfTpImNNUHhK8YWPvDUpsDKHtiKzltSEq7fYLVbaoBueIQh
mXNTK1V8nJNY6pS5VAHpc5ZIL8/Tvm4fnNTW/Z3o6rWgCQHykFtqKHhHVxtCZ2VOZv4vqg5J9ero
JIFGzF7SWrHp1DNOKlt0/ilqCYt66QU/EjA/HvsL8xhJBm0K5kKRF7URZF1A0N6MIFFkr0UEhcQs
C4S8bsfVmH/w3hZ0W+VsR5fN3C2suolv47AjXUGCCtl86f+NfNzVr29qDvJL8qkqd4u+NRBeQjMT
JVdmR6i7o2MxXgQT8o0c4N+eEWnYmzMb5NRX53wTsoSbahqequ/ocoMtQVHGX2kfNqa/KExr6uPL
rtTXMY9ZZUsTNNXGCmDeNRBiiBF6b121bY2bSEhchO1Z8YwvxK0Wx8ZJIme7FyQ1H5EdheWqwtjD
URnXtv7Ih+xuju/L7bR2C9sWreGh5cEXrh5lK/FasEB5o6SvoVgc12MLkeUScdbVcqBsfxw5LNZz
g37vr9kaUirtmMA807HwyWtICz2HwaWxnD12akksxg9bXGYX2z6YBZlJ1/vWwYyViU9yJONtmpIY
Yg+JnV3HGktrnAbMp/WgTtUe5pw3jF6mA7VPpH77hHh63xVRv2v5o5mPSffYO4ZgRRU54ICaZVoe
ONDFNuHYmbDeSP84BGaruO2Bkvtt7M46JUp6ZSqqTUAoNa+vVei6SD/DZnbwWaHliZrzixgpxesa
pgajIH7bMrf/XnHlVjMiFvN7UzsXI/Hr3vHREkpX7IHzd7Hz3stl2De49XEwLRUTMVf5a5MmAeIc
D7gmnkYbHVChf1zBrjVBEZr4MiGh5RdHaLqFPJ/smh1vgfeYdbwZmOS8OBAU4N3uSVQ61LtfPABE
i5v84Mm4A/wWnkeuVz4B8PN24i7dvKTWUVu6yuqdbPPEwD3elXGvZVzobpeupCNB5LvdabEXpr7G
QYiRBqnMft0G7KxaZElXjHRL4rrFdHoziOTt9Ky5danfmE+TX/tc4imVYBHFgvw2XP3d2uutl2ZY
2+NMzcshctPmOkjj1LTyzyrIHB8uB7+X8ZTNiFuECBGgoGkUgcfhrMHataexuUTaY7eZYnd8Foqw
06iP3wsJyIrEvm1AXVpRuGoEYBg64K3HYJb8Uga6DnkY5p0y8fh1C47z2eTBNGOwkXr3kl36jseP
1SV5JtfX0TY/yoItkY6DHhILbQlTiztnIquvf0UY8nPx5gfGNzQn35m/ibK/NAdVuqk+TNPGTBJ0
XLRg0ZEU2ttLbeE+keYSiP523jzkrgpFD5fRYGn3RfV1R3IbB3QhF3vVXDjHmuc0VwvlI6NNHMhC
iIigAm5Q16LkqR7ZI+AG0mOxX0bsk6Dv6Fo4Bj92/ib0GaRIO4FA8i2LElymxONBKgcUwtrasuyg
2DUnuaL1GBubLNFAGGHB+oKD2LwH9tT8nLJGebl5XWP3vxVAknNstW2jpRFv7/+GBs18XZPSPlAl
9AKYnjN5alEznLAk11j8IxQhPid3jfxT/tsodkDcDSmte+djOV77KCLrI//7ZI+HIHhHsVElueWx
WfziQr65F6LQlP7UYRxvBixBuxf1m1J1uzW0aovuh1bNMbac2Lp15WRZnDGqkkZzZRsrarG4bImC
0UnzmSagWTG3cErnC4ePvuLgWS0kIkSjjm1lek72FSRbgCuorK6E8sJApWD5EMSADT+s/GR/iIcc
fKMS03MlBa1cGGLKqtvLD3nYFviLJLuTqW9GCL6NBnAr1UBrmcopE1rc2upkuG+ZTsFOhjt+ePuV
FjHi3DjlCHJ8zwH9Gc6MiymZgFIS2t1Ej3obUxX+C2mx9pNHgnV/UFBUfwzZvMdJv6tkCcV1uGCS
Np8nZY7ePnVIyx1pYk1dgC5A54W/Xa6cw4kl7hJHrg4E8HylgZ/uDUCvaIfUQfvIqbevw9pIAyZ0
LpkJGxfUwUJ9PJ+vbhHsFLNeTixtp9VvCYF6+KSTGLJIUzmX5JorDAO7XLG8vmAaf/okNdtdq1Wf
DZtuY+kNCapCpDTSIHWorKttePDJO9RG2qalZORnHfSBTHmdaW2KLbVeyFVd1B7KD19o0/Vm+A+C
aNMyfQLmqpsuhy5I2SCvBQMZvkndFqII9+bbIvNEL/71plFvsRfPgTcXiklarBgBfEl7GrhomzZy
DrVcviXUV7GfnZEzh6tt5YdiyMbtSWRaRaiA1yeOkBnx1Vkb2ZRsUrnd4GQ+QJOQMFYXt/JnqDKK
cjwftlSI+EKBFkY+dzaoj2aCYLcb2uBIzGhAouTQmh8EfHOAP5O+zKl3x/GYvwa1ksPHFh/2sgC+
39K7EqwO7kEk0D+ICByHkrQa74DUO0mUEteBRWkgdoOjM//0i0b8vFSJXKGAXPwsIPySYBjVvLjb
FFZLjfx7apoX+EInRc07VF3Yqvfm5dnz7HFpDfSRw9xubsl3TQyr0f6Jq/VzfQpMUQsnaDjMTMIW
m7CRhDDq8i/CHhUujL9gtKmcPt18AZNgQEnADSGqjReu2eMdJ9mIaCuo05tC3UkHISmtpytDgWN+
xwMAvkXLfDxNFzyoEizk7EsvorGGZmDAz9zDV//4cPqQoDLnp9uREiFVLinrLWSyIyEspk/J9tGw
Ch9QR3wK3zl5fv//fzXn7CFd1wCmmsSJCvQgdlQlec7FGldPheEH1d5FtSGcuj2PdDD7Tt3npu8a
+aIjRBvYQU9vIbYXRGNcQ4207O/jGA7gEPWe7X0FZEriHBsaJPZbuMTzyvJ8JI2KRzKy9eWu5S0/
jxW4ZfRd4s8sF3ocbYbLpuphvlDkGADomKPZTS9j0si4KcKyKI4wqU/XVQa0XM+CUO8MWIgCSbyD
Rl75cPSkEfEgQqD5CkxDlUB8rkaPXCyhuX5G7RwGpw8wpLVwQTzRipazV9OXdDYkptP26IKdHSnI
6XbwLoBmqjauKPwAjfs2NWIF4lyAcKe+2Ch1hPFwOnF+dO29uiNWZ20TutWpHznZocU0acygBSal
UVmRjeNTdBdZ5bMTuCUtUrP0THcYcqKELSAJ+uNWkkLQqu6qFx78iKFmW3hOcVynpCKwxoP98e7l
7Fb4iEPr0lkKi8zd/XV8va6QkudRPLieJcU3k4w7sP/5TheF/fow43yS0QLk7k3oP0YHvQg/0p5F
drzzyzv4xMGSQb8ajqfV+t0SsaaKId8/bnhxVkey/uUDkdwQgqWIaB1/sTh36aIQNefJlVyaum2D
SV/wBqr2BrPeypdatzLN6eX66FaB6cL0qmc+8vdCbr6GFWLQy6QleftUiG0i+hbaqSx43RTfJp9F
wljLeRKqIgNnbaX5RpqFl6LYpD5JTvuLEH0V5SkINnCC9OSltO/ImzZssagmYgvjleRqoPv9QVOm
LmP4BVNauUIxIBwgGEVOwSs0oITmC8/ztTzqHsVaUSHfjmMPHr4WT5VqzQ71G0wRmTaVGcsVVa7m
hkZxe9MLKKuAo2BZRNcXRZJmBmaEwEMJL/oOBT5z1Pk3czIPaIsL8u6H7/TRO3HL2adHZ686zpoL
WWahMw+qrekXcClmx21I3FV9NjLDy7tQX7aHwNWx56l/n31pcmz/gGmQ0I8ARySbmIPAoIPQYR99
2J3v6RqC5P+ZruiQ1IBpj6JvlhJYpkWMTCGw3ABu9s9RnzItNiyNYFQETRODhgAMntfCErkRpG3X
cqn0A5vzGGIVt5gLESAyNuNZPcpTCDA0duo1T/kKAIWe5HKb2MMu7GmsUQOCFt8gyPAlpbcWrrCI
3sGsLZrTsu2YYjvx5xwUG9azsswBFohQfuhnIAfJHbhk/Nc6eDYwmFhkrnJxC4aeZKijB/U/i0Bz
uY5yATuQtXWfPhqwEzyTJtLGKO0btT9PKgZgoT2VjUIruMVUqxrYiPta9MFKh0kgML+t4l3fZWe9
yvpglYH4evzNWl3f0h/DEiBssBWmExKgWcxN3n2AdN56pjac5hDtpywQN/lycZhTyGFSiefQy20M
1LZGRGj47pvFD1KSLXCMaBT9geZ5d6ck50GlRXOB4yyvQFBo0pjY+VOWZeAo2CixRSHbtFH0nSw3
POV/uoJeGtD9zEqI9WPV3Bxj1sNiy2WoIsyp2N5pkQoIkzrizeX703tiKAhLrMvkR71PNdYXorOI
V+0nWepiVFB7DVqfZRg6/fhGc65JziWpsS32Rz9I7dF3KfbLKw4+qS6IA0/XtT57gfa+hoPy+mjU
6ZxvBuTfQb0SZ0iDdKNj3uXUWA/BGi6QHfbpH50dfrK04c6/j9HVjQ58GsfjHkO6wd12EGQM4tg1
wbLMsSf5F3MPt3ElGRXq0+OqF3WUH1Gy/UDImIKYqQUBR/VelCiuVdrM4dVMOX6+9YRiDzvk1AQV
NGCswLAsD8BPk5SlKkpE1+5T7mVJmCTgRQRupGrMwyMN8YjS5cyF3/eIS045otviHPFGObebU6CT
XsZn45A3XQBhzZOXOwtmyiH+tRVnnCO+1nnXXhrQkpWk4CKVYHM9OZBU3h//xpFC3qh1mXZOxNSS
TVkmL4PWy7O/NugDK5khJAHjcZaYxuHGvO2a0hQPg5trTfG4PCj0EnvSeTBjncOTNih31YURplyd
dEzPpFPxi3xrC914EKu13m6ziAF8W8eFI9cO7umenrfC+WSK5PeW65HZtAlKL9AalMTVw1n5XaCW
vvr7kdgCLtkpsLRca30G1jYC7i2rb/tTeboGbnKIEDc1J02UaTAaW9QYQNhlxZFpi00nEOu8LT6P
WIIeZDmwVGsyntPHUVRBx5awIu424+7GSoz+ga6hEod+UN8uWIBtCEUfXfACifYZU82zjml1stWm
4tidwM3YrgKJcuWZdJFwTBi9h6almY7l5FAM08RzVsxa9fQSeh1CInjhYRKcN1joqqqlPzIc16VB
HQLSRNkFt/L4u7mjXPwkk8oEmIiux5cFo7sGa/n9fIqr2q6k9834g4eaZQzTjpAMebjiQwa+tLh0
0bLcsq4eAfIE5R8UcP1Vdmbx7vqSuK9iGO5/yXW5NQNGMuwSbaT9iP/RAjq9dUjpSZIUOql75K1C
Z4xNbakxZ13vOUw2wTGgUAOMQAjoyw73yMQOIVfewXXR79sZrCRedZywOo6cahsqpkGDEb6alW9E
SZ4fIMsRYIGiPNZmaYhs3g9rzAQ/R9LrN6rWT4J3u12wpqAVollyvPGSAgod3cEq+6R0DVdv9KOn
WhRSGcR1NjuzBUNOqm9Sqq8QWsPBoGlNcO/bgXOV6u0q6NFF8iiABlDqpkXOxWrq2b11x4jiAE4K
MWL3ptJP4rCLzpJxk2LjkR0BEEOpL7Aq5YpmUQg/guaH8DSXgLqJD5Kb5rySu7yeBolsb5zMGqBX
mWeasiFmQPPFOY3xjUlD1iOLq0FsJY4W2pIqWzKgMOcwvSouBdDhA4LsuWg9WDNM+ygxOjqYARa9
NZKo7zfU4lJEedeHLBFpx9+uzaGnNLiojfTITFolrM+/U5hgZMHfGxDSaqJFN7ZrHU+eTj9rnR7M
FUyRaSBmx+RGXSMEFHxl5O2stttzv0g5Li1jrpvrm6LwV8vMBK3o8jdVk0MFt1/d/Ha64Q4qIzrt
ZidmliKL4ZdA5ijFyIP6PPikLipQuknW4F1tXmZDNCz8PuuP4thBat28/l8gEJh1twWbpIZ3RWub
hYvE4VtBuVa+K3floB8rmWSePjdqLfs3XiZ0Bfvo7LC9Fu8b3T5O7QjrwmQOWN6I1DGqIyLU4152
tXqz4k1pwvlyGdyt7l5noHFt9IjCF3873BKbvbyJcQAqa0ecdAeu/QFJpQctY3zwVk9TH7R2YfNT
epNsUbTYDM8YZT+01RkeN9ou8ccV+WU64/0MY60d9IFkf1gyB4q2QIMa+v894UzXdlJzxq7n6U4K
f09gojdF6go9/snzBTWhVAhHQGfwguOIA4d8V7MTKeJ2aMx5+gp1EEPyAKmjMdWO1ZfoGc5Dupz+
EY4BiVL/U1oQpCuzUh1J72FqbUHoMqDdObbT3+F3tTdgUDGwG4pweQFhouITHILl02/r/owOLGmT
kcwKvWYPHIXgoPQdLc6Dw/ExUnDzfyBU4Ao6beCtocBGHmC/Be9jWDWb226RKSOQafGGnfBDLb6Z
hjR073CvW+p384Cxw5e0aVr5VfF/I2uk7lXe00jpCtXPq11vDX0DElGVf385ssq8v/QYCja7UiE3
A64egAuhKgHhCkJN6c6MG1SHhCsrn6xQuB9j5WKL0NTO7ELfpBoOEq725xpnlQiVHK/bCi+pghSd
3NiYYElEuYQA31o3HYMvuTCwL7GnCgKYiT6G4U6JDBqVOpNPHGYG51kOdrVnM9FQg9pBaWE8HzP2
LZ74Odmj+pyNMemFGbG5dkjdJnDqtncvGjgL46umyNzQGm2pL+hK9+PolUC/xy6jS/FdYk+7Dbo4
uqMBjai39KA8XApALiKqxySEJ7f/9uT0Cnv5KLEEtHsQQ64wXVRHjpZ4kBh+k5R/xxn3NMb/zdPr
CVJgz2rPjUSH2t1crkRPZy16a2cnFA9EKuo8sNWwH4K/B9JXDgtB2VNkmEoEQQqn7Aw/FMSgH/FY
M6dcVifxcdqt9+sqiHjL0KzSvdG9vl8LrQ2C2fH4KbkGbX49e3tmrWcc/Ko9Lbl71H6gUIOpJxnR
q2BS7VSUFDYpu95gsTmDZh+xKXtAWtDqBBY0GvF4q1pg3XkU4rCKqwuBMU9IhOXvAupd03ZIhN9f
PGBduNwK5CFBvrYcpN1nfXuHmk9dv4mr7M2lwaZm+AZNqVmi565RRaUoPj4QftGzZjamTyCIeDM/
SPWCebod/1zQeaWG1/AEeVCKB3jlVrKKKHefFCYUIl1higuTlTEtZ7l/e16ymmI/8b3zyiH+BFUU
dm27ugvB1VbeygwLmdw6HMbs/zy/tq3SR/ulOqkni78NaqQnIplPcMLl+le/oGOifuQS1MBFlvqr
p8cojm0zYgAGyQei754+1ZpabhjQWnSxH2eIu6H4k1oue/12KGLL5SGp+ZujHTuB/mDszXqi/kqN
zvyl8J23r5FXmt8Xh1eXHhVfo+fgsthWHMGAxsZel9R1kWSavylr/UsszgZSr59jzZRcyn0zJaTV
zAzwxee5KlqSkhUzWjE3eUFep+UuNKl7/NRvHPIJBnCeLITzIJToYOCK4Tp3Fnq8SIuozGBNWs2/
EA8iqiSHoXAF2oq5f2KsRCv3sdXC560ACacK1+z4I95AWClH70V8BczaFPJs/Jmxw1YdzXUljau4
0uG7ZpLNBQEMIb0YHGlUt/63PDe6F6QfAMosWhB1FM428efuU5xvb4YkKGF/JJXrKbe02H3N8prM
h9G5nM+qncc68yWO8Gpwrjoh0jHOmNpQV0j9HGev6oh6pduRGajFCeyf6L4SUkn7QGAprNv9L/dm
SPxPRpquysSvOiu30MQhw8cYKJhhAOTjaVqNFaRdxzKdUPLOCNyIHckBUrQsokoaTvBvSnRmH4Zk
NXfSXvoHYr74KlHo9ok8iDYkWf8B6mi/BZ5fcsILXAZy3YlXZ+oHu24qp/Dh8A2HITEBOZGr2fiV
qEAI55/1+gWq7hqvT2530m6SSC8hHc2Awo6L49EGSwUsi09rPk2do8UFdwXa6H5Q4Cj8sNrfiubO
RN9hR4RXUPHT33fl5lEVW+kkhxzIlP6ierd+bbk2B+ZR9xqqfuAOHQMMj6C+AeGYNmBXaQUrwvZp
Fi2Gyw3EiGSan8l4Vu4O4QCdDHtqTJTckLhC7ProveOOae1S5ukKlt9Yzo4k2VYX2NN8T8L+Cycr
i85tAri9MpgIEh5U98jRFPuoP0tNuc0w5sR2AoifZLcFrhQYjTcKj3S+cVAKcK9CMZLqlz0cIg3m
jVU+rSMDVYvKDIkgiLocgtm45HH74t0Opo50i3Y4c0luXHvL5Iq0WbpzLAfxB2bhnQHU+j3k/8qW
DF78Rf7Tus1NpfpOkVv//S6i3eXmMAMxKQerV/TkD5tBxIG9LQl5vRoKSFWbmKJX+Cp3qeiVg1Ju
0oAMYUjhdHu3bXBCz3pYUnknm6vYY82LPfyz1SiDMxlFs3TU4DVqkUHujOqX1rL42gPUFUZW+xN/
Ta4Hre7BU0Ab6D/IYN6vnSGXSZ26oqrX74aOuvWONWk5F0XdaQs4zKH9GcK0vuqodiIYRqBbjWsy
prOw5mfcJPXh8zRdqQsRQgdpyOoRizs+Lqxfok2uQW1UUBEEaqtd3wiONvRmnf0Bx+5+hn8rdbsJ
6mr4TCDOYmUCkHUWZYobWUv7WINUwWEAvdfRseeL+yluX+Hy8v1LaOKl5jPWctkWbjh2x8RX6Gkr
ahPPzbikOi8sa2qYEfszrhKXwLBKq+7XxypZHK0ITRRFReIx/2fsbglyLZJA/xVNiAgQmLRGJgJn
XINIlpZ9UntfWDpZxUjJwzPoQmGi4GViRGMFTpdjB6lruj9e1sR2jiFYyCiDNguY+KEYW/VRk9kc
4uzZxxASTIDDdVaY+wo0PYf56TxLDI2ifLlHer+p60Ude9p9MTfLclK645pGioxBLEPE3WiJaTk3
Tw4YSuRSyhHJl6XFsC+lgCL4clgTipbF5RdFfXKtjAwykc0CBWa3b5HWZI489GF6iFsv06qxRnMu
M/6qvwblrrtLL3cLa2xUpfGl0KiX0UBlZUjSO6/9o9rV1jcMms0x6XD452VQZqtvTcfgR/zaW7zT
SqQguPGyICpzvWSjAG1w6Y6Qzy27J2xRjABs16pjIfpfHLM4ScUvjyJekZtUN51k7dPbE6UWzK8I
3NZtI7DBBdmyc+WowrvAPA20Qx6cPYhx06KOA+YS3hBOavkeny1qCY+23AVNrxfWKS2soCh+SPcg
Zxrl/yEvaOfHNtQogFNNCnfVEK5d0bl6TuMNCsrzF2EKsK3G/mxfBv9GBpmvj3xZTuHnNvydtNF6
fTCbq4XeK9kUmdmLyBmafdQyskukM/i2qJBCC8vvgg5UXh0YIwV0G0pK86F3BRY8goFM4S/bn8uA
WRfrv6IWCgVWemcvJpjl8wPReBNm5123dY1n9EGeN8f9e5JVcmL3P66CLB6+8S7zeR4O28mcFqsH
RTTITKXCmeKlXqTvBWe0rfo2cktmD/AaXqMmnR2wGMHvnxrhWbS7oqGW9X2dmSLz5lwaBdt4z92H
EoDgrRDgcD6gq8p6aKsGHbZdS3fSz783IyJ8uLCr2eZwX3i9Jcz7foX3CZNM4ULfieWyRYBADzee
2oxhja0t9IGVO1NrQJJwLnE1gAitHKeKOBGRSBgvDLClIhJrTE00eMeYW4addg5xZjd4ac37Srcj
lY4SWFU/ZKOaQlBqjJZBpGaScXQopVK/JlzGbxC5oxX7kv8vPaVn3vpQwVzkXCYC+prrficpXvX+
7UW3evpQQp92yIhv6Q/gWKSRWWVCkmzffD+P6KdoGKsceTghyIN0ncDv3fHslYVLWubWgt+k7IiA
TWGi6rGCgp0gyIqC9lMlwTANwRHi4wYTcyfjYQtDjehNxOLKvhdeLCmDngpWBLYUwd5E2HLsTaIT
3H/iWHOl5hNheKTrdbeLtrxNzmPO8jLBRsvYVnOtsSiAWYSc8T94mIXGS5kNrsOirAo4xwEkv8Tx
gAO6ZYWAEpChesfSads7SEg2JXIQzRhkYIVHdauuHK9EP8ZwuW0pZMCU/PQQhTOaIAnw0pOMYpWu
Z5lGs8C1VIMc2L0Sh0/O0Tqks+soVwXq/lvSPa1QYqJdFaeGThMy9UexRYuEfDhTfML3/FUc9XPZ
XRHHkDywqZ0FzhRkGSjI8oBRukrmq9/Jf89+ZoFg64UpI79CTLzO331YFz4W1wiSV6pS5okWifpJ
Ng0R7GL+bJWCSLoxlo3dCFyee3KCIbCIHz++FL80YiG8iEWAdvKWrryU2zIHUnUP9y45n/gYE30l
adBC3e9UOw+5OuZlmmFsoZhFfsMdEgh1zt4mIHRgy3rqvtOq3zrrgCNNVr0I9uLSYtMkWnshWnZe
y0nzpuAMV6Z88+VHnEKxy+wagU7by7uh2OtIvSTqCNSPn6D5jtRmsAocqnOddWGHUUUDtCZfCqsL
jGVwLuA3zWpIaQVonrJWxAT6w+TdCy4DDVijEcC4G8f0cFtoECNA2+XxCmW/4Mc01z2NWWFhQSNr
pJeGrBUeePzWgJ2FQyRLaEbhK/WO8LyU/qsboKwealdE8C/UQIbHX8hy5AjjT4R+Dn7gDVpCQaZB
EqpEZxOg8P9JRY7vU90S6MuBmJOhKMk0oXEbqLDKimTjULY6Dts8ReFWA2qtTKpt16+0zRzoypCB
0/IgqDHfCFrLdCKpa8HSLMaMZHT1s3UcninHz0tM/eDr1Fqj/KvVcZxPXvrZ/ACb0ecyVt8V6nI9
OuDYP+MuPQ/A7vsnG1iiyYMaqorDc4viLBKXPYnxDyaZd5cJreLMIgumMcBQ13GNidfDG4enwVJa
A0scGT/Jr18rdw9DTUyxoO4avCPifmRWYQZE+fnICIFHDAH/xEyk3CW+D+ulJYpAQY6G3HBuMc5v
sURh3Zq1ZjpwStGxXqdNFYbMezDVsm5jMc+8LOEBdvyj5ztQwq9ZhGFf8lrw89SOviyehyNhkvir
pL+YIqsTKwTtUMNWyc5Mb5K7eYG3baDgKcHFmFlSFyM8zkjYk8hfvgRvG/c30MGlY+pSHxO59C2V
VSitOwR1gRu+P1VQ+tpTsBz8OV2HyoFw0/ciAh+CSx+8QipU4ZwbWXkSgk80lla6t3QL0Dk1ClSA
z8OuDX3PcFbnnOv4CRZS+vcSc8y+uNxkO++wmsvFO5P6IVtg9fefXWBSyrM1EHTt3TcFXPR0OmNc
tMiZIquBeOoCzyw0XfH1aNLQ/RtDHIQuW5ourMZQcffiUmTqnSRUSiAmzgMcBH7CCQ0G54EDz5Dn
yFR+0GJZhmSbvRAdjnMOoFKbwJ+EEx0ZwHWSK1hVG+hd2XjBKcMeeT+WGmOxlO/3KEKyiZO+B+kv
jUxkjJupvNxFDufyJgHxLd9qL/ulUJSM5a8qezXH4JbNVkjHJ6b08/0/zaozmpXcqaF+XeWDu/ck
cKs7B94SuaqLdxSh+Csf37NOv3sPKr++2DGy4yt8UmcKAwvVGAsefKQ0t6NV9TXywCL3ntpUcnxf
iEXeU13fm754BzKguNRQKP8RRZHx0hgkJtmR1gJIPSWziK1pMBiMo/G8ZeFhpJlXnNeVTxlhubII
CXDBviCgplGdAG5O7JApJHu/Xv6b9TGkppB+uIaq8NrIWHLwp5gZaKKnfWuns007+dqIFFqAG01W
d9dnRilErReR90vjdAjkDh+vxlvKYJ+hV93wUcn+72bPjqzkVhLge1DgMR2EUwKc232tqfRmwOfz
sidDgbe1Z0p1CNnEfxue/5pDfbCEv/etB9C31Vd56U2VGSsAvalTrLPoPLdHZ2JFW0D+N5kN+d5J
hHNyNlfI5GxMMDDbESiUyb11W84LtwWZ+0UipwyED35AbRoCssTwYIvZG+6cYe4Qkm2v24ebiako
oWqHhqbg/zS5DxDS3HzrUUnsng3XrkZfIIfsPRqgO3H3xrGdtFydVKxN0VnlgIsX355PguEzqy2i
HiTBuE3BaoGCm0WlmPG4dvLaaFisoYfJRn9HS6Nt3UjrGYAuuY6bNMOuqXFbkxH8xw7rFnBLJ1Gl
qHwB3VhOgOlE0pf4yiqxDl7sIO/h+kNr1VvHP3TBuQUEr7wsbYJaj72Fl6XuuAwSWQCOK3kSGM+m
7dYc0NjECjS1Wg4MfL2YlAv8zNxcQLqhk/5LYllprQfLiFmWc5GvoLLdi03apHHaLPEUPS7WS9aK
s/Ut7g1/GfizlMuMJOHKJr9CWCvZwSQjCh8FM0/IeRCaf7NUmxi6TB+a9i5mingDL+UjTKqC9tFM
wC06qBV437bgZRSSGayuXtf3n8LVIpWhuPj2LZe12jh68CRFOg1wF6iEeVL43ya0w/yg7ZGxX+y7
KZEe8iliot02gPpaytOfUAbQMyoj4Q8/gNhxWdaRl5rmFnygOwo0Tq8OtOJ9L0w9bD/WtJMo8V09
pQOBiaI6rvyAh20RUSgr6sxyW+iuf+4XOXshKB7XrZGaYQ/bdzKZ8FcD2bLdXFPSTLDWwfcTqJm/
weeYpdYwI9zVSdWq6CWRaPBQOg3i/4GQhPqzKgxbvEzl/hy/jpnXB9NGTj1EuRydTNfv1AQ5xsyU
auy5bgKpyHJfREZLAyNzOV+y0f1CqOfTotxqzJGR9dgviGyvYpqf+OxiUcQWwsNjj3gsgmscleqJ
USQcLQw8+tcFEr7Nq46umTRty6xjT0jrRICsU9/4hW4Ebj5KNwtIkDHewghwZ7wT1kYcPKVRNa4L
zSNUlZqCpWURNYaGuJISzl2t5eHWRMP21a2hkOOg9cjmtahsVTpvAl+DxVPp0ig+GCpi3HTIkc30
IuB7vRFHxDLjx9wihoRwiATW0z+9Ziz9mQrq+t9jW8qA828eUxGGMkKjj+Ak3iGqQkd35TsDqUJ/
V3ciWZqS0LXn/j3h1ddjLiwLrv7dk7T64KmTRcXVp8X2/9MwKtULqYOu0GIfpPCCHGm4OGHluIlX
HnM4yCoum5CqHvRHYjuo6kEtI+wpHsxfH9JwV/+KmZ4OCZN8ftslYsNgYhlTTOxT9iNkRq3LXgod
TcaOlvW7S0zf8Sg9/qNXASUVzS6dIjvXJywIhScjXVCjGvQQZfnynli1zJMRgaD4ZTw1vR7Im9Ks
7TMIVMQxi7rIL7uG7tLBjUJPxinbPVx+6ozOpHg+v72ttn69xDjGmcKP4zsj0cjAFY8rsM8Y38rO
qq1z/Y62jgpIuMWTIwSJY29IDkSfwSqojJd1qJvfM4YLWEsQbcI0cCHK6njZlxKgI23jdNW7r5S1
v1gE2rew8bsZny7NoMF+YTAvjb5UR/aB+iSc62rsMcIoq5pDOaotSTCQ57UjQdDJPCVHgbnswsF+
hXrZaUF9aqJMqnUgc4hTO/FUVTT2G5HrB+HNSjeHNVZodoETvpMSdDauoNHBRQJD73JTwNDZ8YlL
usXQHMO4mn+gpPbEeiN9jwgVPL4YoTHeV4x2wZDAGqW8zpHeZt5zYodxE2bHznrKLwIYfTb2zOPF
HZboeRdvkksD1cartL8TEzPW8B2pSU7RvpYWqOiCSe9zzRT6Q1PrtO7Ifw8jZGbx0Q/ttYek2+Ry
e8kgI/j1PLkm1TwtNqnvnS0kpGbimSqnX7g90NX52v350K/Ql87oyx2nGYAb0/bZi9JOwtDDVKKM
7hzNihkYhICX9MTmYAgz8BgemhCqSX/Z4iNj3X1uCVdO9nIXRFaxyD8MspD3K4lFkWye6QvmsZzd
lYdaTnCZqCgykyMiajq3VjUrCpZ0O0Fv0PHQma5zeE9R8uJchRqsYfRTrBtvVthbE75aXZabK3Fu
b31nxXhMTUlUDckgQCyeZ9Y2yR79DnpbLy5jmlGnUtTO639MADNi4IuWGz6lwlX1orM3GuefMQIh
Sdw2eE4YJaJhyj52bHM9hYFH5aYjCAlKxmX5otzkSNhaT1NlxX0msyIM7qle2Yvu5C4xuxvFIruM
NrzgtzGgz+sXFIcYLmf+k3dDurCS2mebNUFYGfp96HA8afQNKkzNio+yfPQGi6ytlfZt+y8mjp/B
tTxA3YzWpV2UhQ61ASAw6ePBbdvqRWG3Kyz+SkIpr2nn1479qdwVWtnbKrUF+s7ISpfzAoCzhfr4
ATDAmO+1WRrmmOJASXEQuH7sm52KElIoJll/vKaJsTJZ1Et072MmEEzS1kmD0Wwb015jYbtP2GuA
PPZAtweg4yODB6tFFKgmq9WtBtLpAtAxWYwQ9rZkWlZuCfiH9C3pu/GQ6OqMFF6B6p7I7JnSjBY/
LBqJb2KuelwGhccGhxu/AVCmjbVhUY0P0Lk7h6dqR+x8gxEg+YJ5jg4k8fAmZGlZZdMbQVaG/7T1
oS4xdU4fRe4eoht2Qar24GuKCGKY1moxYI8DJcGfRncWmqpLoyhHDjU54V/GczGQ2i1FblDNAJuQ
wGp8GIhrCxwlEAN2uD1jWw4PKdEmrZ2nbyiAQSiXYbJWs0Te3+jYIDCQWGMGiPmEmXZM1Z7sinRE
iEZNL6dN5e5H/XxOZIih8Go/ZzHViJZGz1lbzz3re3x4dlEvrHUtTdV/LaII7jSrPcDrRKu0BO1q
sjAcAGqV2JPBkhNB52qoWPGQu6z/bPpsFwEzUfevWeqUb316Z5iaIxk6sW04KzaSIZywhG0j0aXg
TtR9a6V3gpH90G4doQGHmPe7ShfIxBzA6ux84D4qwZYL50GUqySwo7KqDDptEPX+f+VMU1P8UUch
ef50SuPhQNSflyYETWVnwEPrXDz76/+Z8RL2QrFnoBCp6eeFNsgh/4Q8FdHTO7SnuKcooH5nDnG3
JGx9ZYvXOTq44ISJpeTeNVHdiMKEjsmQUCMEX2q5ZCUKmUCFVPydVymlxb9PrUyq3cvlmajGG8f3
o2aiWW/riQyu9ylkN4pkg+MOy5eDdxBsfAttLJCQUS7mRJt+LpWEYt9W8wg8CD5dh59mL2peDM5m
JWe+MczuboWcaOuj2xDmNtBV2TretlAt4amE28DiOymH83w5iFq1Yzr5DKiSSiJW5F/ER2VZQkSM
5PHZxdxs9SLBBwROD1NpU0Zf5b6xYAp4fLS3zhSjUFsQ4fRK/DhUw+Cb6y80adCvy7hkvGueFgmq
qlZtzhHNBm3pBRC6v1GXrZM1bzzuGpb709yR22dpbe+Rix7NGewTfVA+43jHn9nJy+od9Iu+Ikyc
CyBc8pqTmJVgvnAORyTpnx9wsjONxhyPB4ncPqnBcB4yK+TGFqTq7/te1kdAY6wsjzopaqVDr1Zz
27S2Fv3fE4YY9AxPKfwxrilnMMpJzVv55JGxqn7erZW6me/6JfYB0BPas6aKUw5hGs3qF8AX0A6Q
Wp/6xo+ArwPLtcQgArxR/J141SlvFndfCX6majdlKFI1P2CdB0VtWNW8s0h9zDpAsZfk2HPA2HsQ
58jpDhYhVB5677bSX4PX5uqKaHkMu/yZQawXfEMCdAnp0rUGuint4kk5jgWNzLmFI4kRNioJNcri
BmKuHd13M3E9X2ymgVtAuTDZLqR+if3gh3YP+ZBVG/n26V+KG9xFKXfyTwpNhBIwrLXL+aNZFHOy
hXgyRtS4zCxjVs4HSjuvogKtTwlStPwsEEjL7rotKeAIlo0IJ0FVBVz8uAsivJG7MILbln5z46yx
GrkU0aCgq9jxE5YprtIJdj+X829lJAbvwWyVxmyCzTydCd+nMD/Ya1YHuB0SZX0Iqzw6+76cj266
3rPJPCrvoadKv8JaBa1EjDojJX8XQ6i0FaWsggYh0jSxciNrjZv3mSoRi4S1YfExZJorE3Dzzjku
REoVQkQWYICRqDnOMI09XWgmclGnTvG42UNXKX45iZBRJoluq3NX7pJzTNVJj3tjyGiI8jQIgEac
RGvD0DBs1L0moWhEPJGC7ptjKJ+hXuuBv6WqpckNWfudrZbvTmbABX2EMc1xaupXPdAsoWfpF+f3
snkrTrhwzzlcld7OhZlq5dlenf176iC1qInxUpCcVaw+gXEpMacW3EH5TdwH1wMpeVWwH283oimt
RcOHY4Vg1PAiSYdyVLGhvdajaMhsNKU8WupDscUkYp/tRXkX2N+7lAe+svbFAJfqdB2T1knZZ7qp
ai4SePEW6NMfikwns7cvuMqDCHsUXbLBXY4VA+4yIjcjOkvZKZ1rqgQZRnFHsrGqvkxvDC84rNvA
9JFi3lKc+4PpSSPxXYTnJVgh99h7V7hb9dRpbspZi0dPjGx2B9P7qMyUuoxoXVFwFpf6filoqqng
AirkKgr/z8DRj/cj92Zv48dQDLXnabz+oewHe2QRxTFaMLqXvuHSLXdyLhgSRIkwAtFcZ5vO7sgr
orKFZRSYYCjtUrJ5yhMOIg9CtL9N2q3L6RSNr+WNeK2Bu6CXbAZn2Dwlrsb8hz4U5zvcjynSV38r
+1dRQHwkLBFqQlynYdQ1rCgsCY6LSlfLhgPnidVFTke4azgoWalKEzGglI0ED+hDEofIk0RT9/rO
m38mOK0U/t8hCtW5/4UcPGkDzX61Hv7jbSpOHd+XlxwXxD52qsdDyIuKp9qSD9IbXD9+xXmOgVPi
Z4Wx6sCz/gxK1smCDwHtI9gMqInjJ27OY0zTk0A6yn26ECkmLJE8w6FQLeewa+jAlllrX6F19/Z0
9NOfv1QNRe1MrJ6l0FrwqRgxIER/BDrOaxWj2XsyJh2FRMgw2m+ikk6NgkY/VuSbKX5HMRcZ1V8y
/2savyqNw9vaKsB/SgBokFbz16mJG3yafkRSfjq6KhsJ4bZ7cmYyCDcR/K+VrrU5QzY50MChYQiU
EPP304V1nDeTrsmabhHBLAkLS4T3xMGV+OSWR4eSVhhy/OrphcWaOVrHeYQgOhN8JO0YLcR3FtN2
ioAHTNT0n5qjhfStUaGfB147FcshOCrAMKjO+vGXw/hrz7Jf9AEm4jB/oHmUzNA2n+SsmB0QiShD
vnR4aoZObu475+lxM6POnwHt9/H+opSp/iFXQ5fV+zwExjR9Vaq1zP/yW+iCJ92CnQmC7Q6zg0OK
4MY9EDhWhKzZMF341ZXrop0xFjG2BH+mzPjyRxHtKFfowIQveKHi1mMfqVGSgzHlfHZhUVpK+wOz
H21eY70H7kx08GQJ4P0UVqcq0/flyoWu1WBZdXQmdKPUz5KOtnhqy2i8ZUCjnhgJQsbwNYuOtv7S
OY4ym11QJjcYJ12JGsOlYznFQgLBkxLZVxvNnS0m+qJgYkN1nWUDVDVwrLLP/PseQbhnxhAq+HI8
qEFrF43YKGtspB3g3efOnwqMMX6yErfjK5BsHXBYXgkCKtaCOgmuv0fAkCXUyVaPAuDE8gskc54w
Biitut7EtegQfWBZN7Kvjv4ZiSNwGyG+WI6REa8ISBGDrjSQrrJ4yzxRaJEJLoypl//gDUASaWvJ
df2wksL8ZAKLLeGZ46ottPZD095ldUE5sUJfgVPgMMEA97/CwaIlOe8BLkK4Ckt5RCV0hsaFiMyT
F3DkXLrNBHMyagd8i22OUn29Z/P1ZDXdTkqWA1X5FBL50A/BKUKacPgyZ1d+bPWLite6bvf12e6l
hD3koGgpFYpaMV72a+n/cVXYx2ywj6A50vXFlw9YyL5rG2cVEcpaY2VWi+FKns0ii1/nYlJ07dOi
7Lqfjn9bhd85QGU7URtO5od7M3I65Bq4MedeN7aQ6zycLnG0iyOUYCMcE2bPtts5iUPTAk1N1rnd
WuPJsM3H7Ln0AdmnfQ1UcYxua5/A13wHofKUbVIrzQjr0JYoEn+xgXY+68LSt/jyrIl1byQBOsko
CLERRuHks1flRduxKom3C/cxcQg9nwVaf17AyWbQGL8inC8WAFp0lUvqXhMJPxFEmOABZOpIVfpf
6o3T6GbGVSQUsdyde0G4+soNs/TSZ84XbE0CERG9hRpNDx79xPPZKzxi6XvqcK6EBaYjeeM0fwLN
9I1S7m8M2OVgpa+g+YmTOk5wOfDqFJfyBEvLMjnPEiIbv4GLlQZqg4QWmRe2HAODLNgvzrItD/dN
YHLCiefZPGd+TlYeZrNZtjZjR8dm31KNkorh92EH308t+N9YFUEBucGMKp+pVWy0OnWdmmNQAf+M
oqC+lO9IP7eIMedayldr65DveS9qsPAVFpcT28JVR85oPBgX3d7b6qFcNgfRHYFYP2WO1xAEe7aG
H3lbqEcyVaKwFGAM7ICfTw12ngbRjX/czfdL9c6C/aqH6q6Np2BtBqhNr/vIAWCpVjsghWB9Axlh
nstSxe+gloMhA4PkhPLX7j+HPYduyUn34BF1QouJjXl1H8BFgzqxdh9E5+/hvryc19KrbkpfD5Ge
+76wuoDuhOrcx4BOcV4gAHJ34eip9R3fzj1/p5mvb/KCl8B/6aL/E9CDe/nQ/370jCCZK1cssGJO
8iYUB9XL5EUblAJlKA4fMY7Jb+facc7A3i/48PoB09xewgYtrLkaAGjlPRPlvWw9KcOSiudUys0W
C/1/XFKz3JUNwyIyyCUQsWrqwgVjO851zluvY8+S30L+tI51jdOAzcnTaE10h926d1M26ULAYAB6
Qaha04x3kZqDPl0dA4C2EmX0H6RboaZJoR80WydXDIfpY5iISs2n0hQKkENtda6XoUmCSPDR67aK
8BsuFIexCblyM5rEbcz6qd0AfyMQPKdpVXFqQtuz9rkRrA/FfdvhdUJxTiRT1XVQNlB0beWgqSRv
IoHaJfez7/t0kjuSX+IjyJxZCEYdShvRLcfYsxAdL6bIiec5L9WWFIaRtisMQRpSG/tO6zxyOHXN
9KyhhYYlDEAhO4qjhajunaiusHbdhv2OXL6o1ibfkZ0/jk9E27+j/DyQxhKwBZ1QTxo+uYZPl6WY
t5Y2Wfnk3X3lUFeAJ0CzbhnI7g3WB4SM8Cbbzb3W4llqKDQmYsbzeUtzJPq3zwCu31ZZ+F66CuL3
s9Sv6vrLcqPzaS7I1XJij7i/aZDR+uNScPECwu3fcwlxPmbTH7AKLfnU6BbiQdDDULxf99E7EXbZ
+os8X7dGQZjAApsh+/5pscDVXCsrrILGbvI2kXILIJASv6Hc9UbhhR6qFThX86echbzCkrKWLfAw
ds1mA/xw36TNeUpaMFsKQGeBM8iveVlC4kicXVQSHapWVv1zZojB5O/l6JT5vdKYfpp8uv9ZJN5j
5Pdjexm9YhfAjVGyU75URgBMvnjMr89PF6TLmsPW+POBCMjuxxBN6HnAVhGX3JHqt4IWKuJxYdD1
etG+fBRVDkCWa8ojw975UbiFzTRiNgtnR/qjaE/ORZDhT6BBw0NHLuHwtNK1VWi+77QVFhfx2Ziz
qPB64/7bDjxOf7bXbN9fsTYzqLrMcDzq4u44xSgttxvZxeRV8WHazJfUG2qTOkNKWSlADhzPEEmg
sAe+9IOk6R9jTM3rHarrcshqIzBOkgfiDcMOWChUORg+CWhEH5/ENzcfRtxVoAN0k0k0gpzOc+aV
tfhZBI/T/aW/+scWnn/c8WAs8WyBruNziPYwkNDtDYE/R/38lRvkmLaq4w5iZc4ayivdaPTfAOdf
ImPIdn8QPik5zRXtLnwbZDwImu2hOcN2E486POzdSUk7y6hHjm25AT7QA9RBoEYs7YN60Tt+incB
dZbuB376Qo/VZ1Mwfp9xDG2KaKFYPC+n59xyjO29fpnmekLrggNK9PAUCFt5ct8z7BAcGtLk3mX2
EYcNZxcAOODEXwLiapjmdJM11K1PUQpxRe6sD8jQALr/VqrJpt8iRy8DJodvYri9j6rsFheaI14/
Nr2dl59P201toX3U1pAeFveGPL9xAmOfp2Wzy9v/WKbWeqJgVciKYUe7w5sjVeFYePRhtPNPitCj
K7Va2DQoPsxSXZAyxBheSodnV0wNnmzoQzjCnYmVCctPbG8DM1f+Sg1rUFl+8ixFBqeG8ppNbpa/
KN6UHmaZKDX3hiYNrUMVrvjX/w3rnDzmdjD2PpFoiFVsY/9tdcHh8YYWGmGFeWsoR7axibrSF+hc
JoMyeMDmarVnvedwU11wH4zpIpnAd/gRMyoAEWNbMUgHLHrUXPpcoCGQd1L5ddo9z6FOOKev/23b
YwkFJY3TpbLGXb44lCER/irg3BdXMzv9r3XaVRDbimuZgZD7yGKE5CNIFrZE1w0td4VvONXcn7mW
CGG8LmioB3Vvbg+1d7YxBAkh0VlItHCOIM39Aj/g9ApnvU4iEVJi7gKJQy/GkajGMzUDPgdErEZq
k3mvzNkkAgMA1ZQf2zs/LSXYWv3XnOq+K+E51I430Mc0NOxShO7srAWTg39dn9iyBEeijtEnPHW4
BiK+ylPz2uwgjoq7pbES90AIyC6Wz7RWLzBXDSXLBXBaKV4ElckfWXAphxu3fdyoXNQgj6xxrP3L
fEjgd434TyRWBe6aGuwYy+9ArhlREf6tR3rlQblUvButajRwNcSAmYldbXiMxYszBSvfH6qGmhTT
gvibv8jF0TM2/ty1qt0TEeLA2lp2tQqNuFiJwsg/FThmEYCglVV+6MYGYvgIkyfxbwFIaEf0hR3u
oL//4qG2JtRbhs0G5PNQw3esLePfGdDPyLa5H/AWpNlDJwo0F+7PniFm8te8kp2IrmtcR+XEoYHl
dqOYC9xxS/dxQVKSJES77hRtazSpdUYpNxAQBdLEk8K8pCZI9sasJVc9MxaoOuFZbGTbpQWhF2Xz
oozucSCm+u1ipHRmb+Pcz3G+9zlSUM2JpsC171PSJo7qYYBLuq2zYv25hZ+raBrtEqpD9IREbIW9
4arAfilP/7Ufx5i3Cm+LdmFwRTtb+JSDM/ONU0DRFE+Cofs89WbmPnWRx6m7Tu+k11Z4+U4pd7dt
aBqfKjBWq4Vw8MRozSlQVzk7Wo4eXC5owwXC9wfzTm4ZgmDBHWhxOiw2EsdighiUV+4/n3Nc2aSH
UJmccne3JGjZM23jH+SkM22sob2z2HGaeV6By46HjCNUqhayiJGWvOiDymrXgq3G4NbpXu/KYR90
9OgoWAvGcOPZo9m/kbu/4utLwWMMZn1evFhFf1DdXEkFshQn+4ccXsTd1u5ney6X4uV61YFV0jZf
qL/Le8Zc11X1OF7gXP+R6jEzLmaoj2Q7MvitagjfW8lL9l3TkEg4Ske+cgUdq4Vy6hdTAVRgzGpj
O5x+IsQjmcVNWVAj2q1BfE/7kB9o4cEEOm/XyvZ+tof15zsmXNnQ9Ta63q/XkcgzmH+NamnJ0N+l
hsBLXBtzykGzCnY3AjtfH6xI37qLPYwY5+Q9Y4KeI6SG6N2CzF9mEq82gp0lHHk+W97SZYbkKd70
8tS79mLILHVpjuyFiMXvuMcPfQSSe8Vzkk/UYAbQ0vWnP+zZ7bf7Lv01kvm/d5oRpraI33vwH5AS
i5wo7inXChXGfHGm/taGBzwNeHkRGVUDPzvTWmfESP59TeYZfrB+ACxzoo8Sy9uQ7NMal6YOqLTi
6ujkhlPytTcZWwlYQKM6D/zlf62COUd4ZXxfaoOwyBp76LoyzMlZCvENlwoct6duBhanGpkF/ppP
uKKZ3TMgcZML645Rur+2j4uDiek9RMYzz44iuwcP62+HCiJFMPSn4I9nkumipUORGHsABvy180wr
EpNJzgp28eJONRhybwR7CG6N8WR9Bdu4Uf7pTf0S/ju91dkNiO8flAksTvXRmfWJ2FQ6VpaB++dB
323gUAt7j+H0yArvuVrLKcHsCoRnsxSZQbMCtZ60e22oBfLFlKifydRUsCcmGck+ajBU6pjMktMz
ayTFEZq4ffSYF+nPewDEO9sVzTgYQT5Zaq99+wfGX4b2Dlj9pOZyzmrqnJA84Ewtopx8JO2hGmsQ
Yp1JhfoGuFWPhB5PDyo3p18FMuwkTT1Xb/zMqQfqqJB3BqoRgvZW/cY+SWhFSHN1EnKndLOCLjYf
pJZte5SDd0dmHbqWAUUI/ZoXFGW9iFfLBEW85Ge2TpYIv2Z1K7cRkEco2S+Rp0/uPJK/czpfQ1jc
CfJipE+IStzvQbtdyY3G/c0h00Jkk650aiNuXKDZxNLBI/DO+fbOpdtrEHhfX2sdWnGBd4Cg4kzB
PUonDu+sxANXZS0PDaZQ1wXdk2HHdS614u15k8yMEjA8ArSqfKysbJMXVTkA+7909Sb+VZmcMqwy
AkzQ3vF4ArlGL+HLnI3Z6jZO9uoQ4BGjSAJhydrawU7QNQk71Psfb4VI4Tfjc5zcHZBQcP9F692w
s7mDoXg0GpTlZLZrWF+tI3rDY27ipJEEPfrORwtP5l5j/soT9ozLoIU+slcaqhT15Mz60F72jNAF
/6CeIQNPzUaz0aYGxH2+dP/SdkWowh+/R0d6lirfZbtxggJ7BJzYfrjrOeF7qUoTbzFNXySxCjrC
1B+vMUezPzYB9ryyZv1fVJxR9Z0gTDPnV2joqRlHIHKY8cH7FhEkg02F/ibs7qKkl6dlYRi2Ic3E
Fzo74jsfa91YXGWGUwYSzOcPBc56QiIAAFKAAmMycQYs5cMyukZgTrXdSppl5pxEwp4Xt69Dtx/j
m59MXxoLfRM+ZfyBsx5et42/edhPHp/mURxLuw0o6K1VBlxghTvJEJA5kWhaG5oXzJLq7A0aJCQl
221AiXccFCVHpmwUyyIfo1Su1wv++fKiKkzeO8b03OSaiRUfHdELKt6ZU5I5nwsvxZ8F7TiCpM0z
Xm6ZLzcMMo0IV7x4NhzM/8BJyvXRrvrhE6XsOoJfaEpfg7bqpfWhKOSRSl6ZnoLE7w0QIlOzlRIb
1enw+orSPVAJpyt0rt+V0DSGxCZJQIDffn9zk/+qWLP4W4UDm8vSKblaCujYBT4Q+R0xAvgG1x3B
+ubdJ2GmLSrHW+j4nzreHgENvbxedXgmZrEx/mVdFu6Uy8DWwl5yUazPsv3MCmNuQNf619s9FwOF
VI/cEobmHS1Pda2AcMY86g3gcIV73Xeo3ANrWpfToJb49QWXqR0iALphKwdaOf9NrmpG3uARVVZt
edkt8bhBk2CaHCOyRZJkcCFTfKDxc3HrOUO0sfzoX0DGfu1FfiKl90ZUMSV3mvnPZEs9oKP0u/AA
cZ+9AOCC2FMD/AhInon9sw707tAn61aF1/2JcysvmBlSQw0Ey21/9vio/ifD/Ldv8ujkvsqzuv71
fUINfb8TBcrhojW0B6l2Dqte7JFiCMQ5apW3GVoQiexCzYd+E4EfDX0k7RM5fZRRW8neH2lY5maw
apW5w1ftLWz2gSUuBIkeCk0V7teaBO4ObSaWTggM7qyL9SjfwBztgvBxDhXQ/7SbwjHi4XuUZk0K
OI6F57uioLERySSyqdUrStrti/4RlVIDK8VO/5YE5FJSe8z99G3qgaYRZ67iD5s2C2SA1P3S7J0l
1GF4grTvmY2kzWCqU4fVQpIslaLc60EB8vqPGL8f1i0p5U7mPNjnSiVkhFFi0q77aFRA5DNdyaPS
C4tKbMscqertLwzVMrbqChVGHUXOCQKVx1JSIFB9NXBrn96FEys/PdQx8SEl6BomJ+tUS0BILXkZ
qQKujZ7POi3FwZsaZrVy7g8TjWuHw2pzSrWoK7nLpD8amPnvTIdLA4AQckDLKHb+C/k3+8BqIKYl
FrCCmSD3eKtyW05ehIZAsQC/AHMHw1OoqxeHPY94vL2DIh7VsVEUQu+VOs9KG6GbCYqSA7ZF6Dhd
E7RvxkeXUIj5yUmP2mIBY8lAXI86M3sro0IRh9zzdmHJeGjidiqpWHPmfMNVFRQaCDmKoZJOZful
jlvfJCTjU1PYFwFA3e6DXCHIc8QRZbsXmP44+rAEkIDqcgN7CdS2HTGtvOtLx8nn+LUK2rAKwTah
Yh/PZmZsefxDJXdV1a9FGdYOnXDMAZJdQLWiquAdzjPRsZNPLZiKChctIIHZzekwsToZ0rLJHn4U
Z6OacizLjjBo6pW9VWbH1O7hh7a/HeuWuIcASjNK485DGJDU0rfcFyOh7FRu6ig4qPqzQP47Nzkv
sPWHWfiJPngeOgDJtrw0O06BwijwrhR4PWXe2qJ951wqWpuQGqaOX+mO4cUzDgHPuyXd3aO+q6b6
PuUtM0BJAMY/vjcLsrXmtPQfqx55KwMCwoXVMybWRAIWBpOtSu6/U2GT7/aNkWclSkXaLkaguOSf
BNLCbip3SrEVjJkh5AQvx3YXZEMNf285SMCU0dSpHvxqj4g1PhYe/l0lmXCayTUtguqXvDjJaHN4
IwFLqu2BZZoDq/p53vhekKA7XvjwtFEVEBhhjJLcSsrOmHqWQQ+x7sYKmIGZ5YwfBXbmfhXIV0vb
vDgdvlBhILJdlfqY+3MM3yI64Zsn/T82BVcXPiz0vLduUaTn9pDqpIYyB7Ji4Z3cyHClPHSKdDox
L5FBpdS0VKyXMBkmh3p7gtxlFahAyyOe6j1+3K1UhXxvU94KI6YYUS1W9a56SuU7YGuvYbJ9JVob
2I428/TAfPg53dAxGBbfENt/9j3lEckzJfee7fssEi6usg1cBA2iFhPC1QMhe4G0wi/N1LyBr8ze
08pmtyStyBW1NU0T2pkrEqWFHUM6p05sh6FlyoN4QGXvfFw2XSbJrahy6FQgsNf4W2r/AiX8Gxnk
HQHPMIaB5AV5K2OqjmuJzHJNzJCTRCchdDpxliOuzPA7AC2cCm1azvimA6TvUZR5KCp2emD6kNol
jku/o80jvDE01+I3HAjuZf+Yixk1UzBOsdG7NkMtFYoqbp4l9UXaParpAzQyrJGQddS9rNxGPBck
1dhLj+v29xhW1OjWlYcJGnUJZ2Y6HvEhENxmohgH4Ng4DFR5AFay8oMEaWgQv43K3xPcWonHsytG
9xK18uIwlAVjTjc3huHgWjRycA5HbsWI74LoAJ599J6Ep2Q6UvnACHukLKNMbXy8ijkvMZ5uYt43
tOIZiCLmI12lj2eOKt7gB41hfh+EKc812NxXWc3yw8mUOv0ME0euG/t2K+DMVuJauYas6kgHlTHo
fuIyA7eDfR+iROSlSukQiU9svrIdxsIBX/SnL91bPQX879nOS3DxD08ilIPnGpwlIpXjdYJplAT+
iY318WtgJuXycfayTUsOj7XJQDk04RmasCThGf7qmcRjueldHwpDajz114SUsFDxScyYaMOpSckh
6jrD4LJTBbm/3psOaDdA00n97ys2hm37lS/Y4V61BrwF2RUnGyuCYdNyKanWetRZ8SjPrbjrqq2v
kK7c6Mf2HYkjsCcefKFT3YJGwV+gUDbPQtfJFn3+PCXRE6o55+l/DwEQTAZoOUCeAsvtGRxjFO/d
5zvx3mT5VUBR7uLRG+7h87MwxzO7r67unKub/LhaeWZPnncPJD96NsEWzy0fVekC9CIZ6h5OJVlp
S3kiH59xFaDR7lk6WhoI1rezhuysV6y8QLrj84cnPMKgK8gW2HwYUBGr06oe9fBOKFfmqL9LNNVm
N5Xf5Xwb9xhp6Wj2/7ARsorAlP/M7QXXmm/h2EZyn4c4KL1AUhsYF9gIRQzKLtMx7sI0LA1STvTb
7qW4sCFVqRzm/hlmJTPHR8Cv6OAXQl1tZ22RZ+Lg3dF1/JM1YlFaFjp6rHfp1joUuBek0S5IYsjR
P6nuX/VkH4bfpIzaTyGJcsUBtPfMn4BQl4/rCsPiseLEVQ9SF1aEfXN0xminPRj0DF19jSFzKKNS
DOV8itwlJoSRsLTcV5Qf8giTsc/BUUiPCwoW/OxX304wGn5G71FJewf6dLExSmQGCftnwVWjDmgp
8YdcLyN8UnOo0hqfR705wIQwHlgpfbUbXdW3g7OjHX0nsXV0aWF9opXFux3EfIL44B2desULS5TB
rcbrI9q+pu8JB9vU3qeda3uE+/SThZocWPjmoPAi+D9NdCnkZWtkKH6c2k2v4owCMytPWHRaZwn7
Vg7PbElQpA5JcylYY4MHHGGsM7u3pozTnd8eXngwb1QDPb4zai5poVJm+IfmcQIq96BpIbnbsys/
p5IxMTeqzjcigPSN/bt8wBrbyEsiZNeI3EhuG11E1/ICDfVJFou8KNozRLvtZw4RmU55KafmUfgJ
93uF0h4obcf1+o2o19HAZg6OhsAiiR7lrLZcrKMgMNd7M06Ljhpfb0T/FQqztNLelwdooH9AxSkU
J5hEwz/yj+VFI/JgHgM+khNlJ3cZf408U3aElEzONF51EtzMx2J8Maa30hm0bnimTbVBKGBTCiK4
R6l5qNZIbUVlfUmM5UjRVsOdc0tN6gFk90h+DeHONlWj2lWNX3s8LyhdVz02fHoDCvPLVLP5/b2R
WhIz5NHRq2uSNcCWLQUKWdBukr1E4DXiUDUayL7y6XCtuXj/n0SXZ/wfHdz1sVxt0+kNidgDzfie
tvsF8uP+KDUPz+ye8vVj6VBmathwI47Hz9rjnMMFLrb20ZkxiMn0+azmfupe6FMM3I12Uw0sTPhX
9s3O8LMaRx2iYKhyKZWgK4guZrsQqldUTJk3Gs5TU/jvBw3EHKf+SGddia2LT6iFwyWZU1DpP2rD
zgpM63FQyTvlbjWnNaMfvpqpzt1UXflhmJrUL9HUkILgyLNXxH1gu9j7XUsCvrgy2tRZZX62oMtz
IhD4mtkVX73AoiDUSZuby2/P8QdO+CmQUldWfacyqmikP1CWcHtt6jjUT4An8dVxOj64dLTsz79S
KX9k7oV5wSMbi0YR/aasKG/+cLXF/cizvfBao75HFF7j8FFLejEAz+zFEtIqKELjBkg9SxCuuZqX
Im99bENRMUwRA6j07ayey0pqEXl/y+0zzXB87t2uUsoWDv69o+NhfS4fq+ka+Um4byOg5EQ2I5i7
Ut+Kxlsm7ZrcartBoNFjnaFuzHYTaEGd26JtWG/Rbx7ie8zyley17oJ6yUzrltKANdQgHpz1MSWV
1+sfrRRr5hKh2JoW/eKonSiDgqijVTCQopLz9VP6lfwbGn054E4EiBPrgQqVvFqrPetGx2YVVLbE
tqKPz2LTjjU/D/ln3bBa9f0BsGtyCmhngPESfnTzEpPxciVyvWtVzU81R3TuZCikt5/GbJNz29Ql
qxF4aYp05ro0byO03Wf0Acc8IWYjaRHpH3U3FsOvkz9iNVn3SNWNkG2fAF9ks7oQdYt8YkexZqS0
p/YhPnfUbUbwoaT6TnGfc3t2xrm4kn861JEFWBbCzzM4iK1kZb9rZLeJxbECOtfV8ziFrEyv4fwg
tvf4PZHQIAgtwVa3t8Xq0PBOC8sDUKprH/sxM++kTR+r6TOXzXSWpIfzRWvRTr9tu8n4BSNXoI8h
C1nSIpIyaD5HHPGf1EQf/OAh0uLvMEhdtPLEzNTRXXc1cmgERS//bzqjcqklM+0av7U/4mzgttay
ENBAk+RjR8P2qtwy5BIJiAkgqxvnUEgb8FeYXpZzw0TEw2U0zt8enIkAE9ixYskngIc48hAvi4cm
WMGAtjEiqDmOE9LcOqDZd4bMFJteVtP5LwnrAORz0GcquyWYbEbzULO7EMsgOn0qjCwUMpZYMunM
cPKqMFjxz37qqmmzDKHWSsl64H1LLUYN6ooHm1cUtM8blndjF/V8Gzz2oadanWVCmq9tlO/EFUFl
zi321pQrcvJb3VqeyIie4Y+wCahd1MWg8MsdqfXJVx76ggEg5t8ubkgyo0xtTKiaJppfLsVXYtU0
unpa8AvpdmePLbRWi/WqbnsMTFCTqzpYf0fhQ9YlRwnecWMl5tH/Jlt92CMW+5bXD4Aa597j+2P1
uVtfC+7MdOaN+D9hEQ1X1RkU2XzOLdhAWH5fSTP1NrxeUyfO/561kjS4fg11gBhM69B3QhNjw8jo
Fth5PtTnlP6QntIpuwI6UXdqhURpKtQSgcZ6vyqZQPw351/CmRQZe4le2l28BCIyJrqegtXo6MXo
fosEAIIF8DY3HKHiLbKhheC+xxV19Bwf1b9d5fo/z9hNRadQwMoVBnD9EAcGjUkucV+qkMiwGZ42
SyFyzoGktfaDpbAh4nbI50rut90ItTN5eDko21BIiJ4kj781Pyf66hwymzcwBLK4klsSTgYosyvP
9TR8t+Pgmnha6NBlUHis7FTq8hz+zqULcQRgxsja7j+4dvL9QYjpSscRgK3d7je7kDgjGeTArblf
ro4wUPq/9LV/vcKbVbY6G0v9g5rMBmwo8lQP4XYsO1AvKL4FqhWQA9vILtJN337M/T1ZMMDsrbpy
IQS0sb8RnK9nS/D0hhlZvRJdtFwBdSZgMIZCbL0qxcX341VJjM/e7ONm1BBf4T0J0WEmHv3XN7jH
3T1cpAIW8PunZhgGls7/N4IM4XpkcNvcN3eeLZdp9n5H/i8gRxIrHGQQwq6GkCZHCAn5bp5ByT13
i03yjLbICpxAXBTHYNcvQk24LoY7RWSj5kEOuCOCoHBuD9jhE1hIagYvmbogYtlhV4XSF/7RwnDn
FVrKX3zXjV1kU2MJMlR5jcrC2QvXztHMPwV2EglVreddi/jTcqlou/Orco5euAUKDmfD7ECPsOW3
8mXVTsqT7FBaeL8FSoOO0jfslT/ZdARCg8xEtZaRUEO8ePsM2HtAWt34qMFynyUEIFoBD6EERAEe
MsvhI1aHA57eGvI7JjlaBpY8p1gyTf9QuGu/9hHRhCnA0gybjFQq0Hey146h0niIKiohmN1HD0LG
Nfif+8rhUhlcn/0+U02IS4mBDBNqD6z0P1LNakfYrO0Emt6lVseLrIflFTNbQPARlPPH1+kgxK4p
dZ2qBV+v126ZktNOGBkJ/3tLCgnNHu3cV7d+f/+Cm/6hh7W27cCvkbPD6whn8Rxs3GhOhKAtuUyE
LOwEOvcYuvYgGtkO7cYRuTgY7pl6ryEbquD20N+CJ5WF93VyZyVcGq7xC5tDf6FdJRSFJTmb6DoF
x3XGrdTwBIAXaF/KuW7Z8HglTdt/Qq+dxF6YBGRUBPgiiVWkIgCYL6wenUdwThsG3+xe2E6+Vdm6
19Ytmye6lq1Wn67luN3hkaeogT/uZ5O9GS/JFrHY42W7guvWEWwlqr2979cHlak4Qwua5DmHTl8D
b0FlQDPXXv0ByqcsdNyojVECCGRfMepkMH+Ot3e05hkjrvtbPhVXG4o3CuQqhqVy/0EYiWzKishZ
EjI4xizC5vbRLT4j3LrOrIawNxVaY2i9zWp5VO4KJGY1N30TGlz0fZ5oGaDmpEYISi9pNJDFZbPc
U7/O+ISTosx8jiEwPZPiRBckzyqcHSepmE4zCz+C9LwkTGK2IFdIuCbaddEWMgDa84fgRFacRXGs
9A5i9b7/p6bNbd3n9RdSbSM4T75XZfOOC3dokFa+VDXRCjRkRfUt+6/x+DYxhHPExLttzURfY0g0
JN06YtaLOZEAOExkiwDw0SkJhtTGTqqD4UL/u64aKOcWQw8IOfEPLgWnqM9OlP17lOXHNIVBexTh
g5L2sXIkc9uyWOarGXQd9iH/2vtKH8cDCda2zzZE30rkC+Yz19sPfkBrfPPoo5vSklL+u/UGsug6
H2WX3vqdLT0JyyCHDw5H3tUgxGD4nrnSqGQ7onMlRrpX5cTZRmPneQqVS7dr0eY1sjbLpEuO2SjF
W4C7fRCLbEDwP0MHOigOR+PZJmiccjYWTl1FQc4u1jHDRBDeOwUiBh2OaikK26pCwpxChSj9uhW9
HtRFbvDDLQNkWBkdMSIsuGWaTG3salbRy5nRrdq13pZsyBkGhwM1WlqxyNz6Bo9I1iSFMDW747B9
DMdjFfeJtFLOuUonsv7Ilx0pFAIeCqWene5QyT9EhLUqKrNvIEYqB5ksWVtWc41x+4oD8vwT3pk8
fe9hpOvVSQjh9ECPdZwKguav0+VJdxIhouYeUOEXVBwuETva8iDGs3hY1lxecrX5vXuPiamXxkUw
pQ5Lcy+oEC8Nk/SZQj3PUftNglLF5dwuPm0Uosx+g7wd4hZGMsd9N1FZSQ/KJI04srZK7bIjyFzB
iiqVtPYa11I2im8PB4bmSoziy0NHsSn/1p9FsUUfswMEWCkHKL3JSsWPtLWpnT38dIWrUpyjM9WS
lWIar+cWewbiNH23Eyckhv/cY1JLGaojlQIKHd+hqrouCA0k4Y5F/BoFinxTxKShC/FaU2rQ+naq
lrTxSkoMHfqsrRoZuuEoI0A0aIsqFf4EJSL0gVcL9eg2Ow0uJ+Ti004Jvb+a0BiHnx1jCPDCyE7T
RBLm1hFGszUrdWm82J8sZ8GmDmaqaqax/bkQMGJqji/D548lfbMSsglqoImrGksavtkd42A/9OFx
SHBiXgEW2Y/7JfRMCmSGvDzhJQewjhh9OexfK5IGMuGdmCrOPWoaWJ0BBEq6MyYixEhqtpP8cgKz
eyDnw2ixlX5Z3BAA6uhFqT9C6i5XHoHYt+JgI1rmCsMC39yrqFPABK7jyB+3VUTn/rXjKWtYEH9Y
86+gHNbzA6kyFUNOY/aVWV0pqLQiDVLgEDY2gkNGKeBfBshcmdPFX/fv9Pbz/C4PKxwugJXLfzhp
EXZ+9Tqj+yrNH2sy80dN+xPsHRUwmGBsZETfxJnMPszVzr3lGI9UOUz8rmJKVMPAE+1nz0rpQd01
W83Ce9Vp9+L7yFppF2H8NnNfHaWwgfAIredwkv6jth0/KcA8MGDVbnG2t2/gE1BUN7UxKV6XhqyR
oyFNr1ls87L044yXBeM5f0CuLxQ7DqUHY+kGDP2s4uwxG6nbgESRtZ9lOeiPhUUVeA0xT4LC63Ig
yITcgXkt3rBjRI4YHuKZJFvBq2PfERByUGhTm1G5On5re263W6tO3KL3vwYv26P5qdIAKDBO8nE4
ZLZkRY638n6ZNoiMYVdBGrlnOke9B8JqsnAUEzD6CgAqJXTlWan84i9jqgbhKGMMIU+GqALswnpt
Crwec3YJFMp6AzN2QQGwXVBebTLG6oNawbd+sz/1yPw31j7njEkAZN1RCJpMMxZEbAwJwAHgBbKH
xEsA/23Y5p8QlFc8ER1LOsDsT6N42nngcVk337x3uWs25W4HdK66ftZ8CQsm8HnKKYN/z+raVxWq
YVd+i+m7hcvt87MVV5At4G8OBm3iY4QxTWDw91oXXlHuVX9i3vECCR8BYv8ZdlOMFVEA5kbeGWto
9CjEABELf7IhFjQCNSwvvM1dPyoDpXwj46H0sGo+zhvMOWc/Hh3sYxX83WPyzF3E2xBX2dK+2hPC
Z17RMiaYz4dQY+jvCiszKUUGrNSzm3BZm/i8g2cXUz6cOx4lSYqOYzpTxhHCurnX3Au6EZpI8JxB
O6ZsgYxMlRMcyut2Jaqz6kalP3BV77mdWGUU/cWdgmsCfdWp8NLnP6wDP7tluGOMyOOkUH/qdOyQ
aO3wU9tCM8gwAqwBn4iwPalBf10PKd2AwKt76tl1MyZefOsegmEppfHTjw9RpxanxAk5WXew/gfM
cx1/VRqFJrKZG0kW7Oson8QZO1rwIxV9Hb3dCXFf6DuIT+4ijj/DxsAH4BEhy7a65eRTtrfHKVa1
DnZlstnSqStNfwncKJNA6vHGPkjCIXpWksOQGQEAanmEUSQHNj2by46jvKSdaQiumgVBzAKvG7+I
AeKXofIECC5nCCTXQRsOFdh98UAb2Cdt/r3bA7Xmcds+KfvRWXK6ZXac91VyBTEnM20rIBEcxeYC
4OZRhrZkSF6jrki+cUo/OsyzSvMgIZf59zdpp9DvXqYvffduI2Yt7ITKodjXS55U0TzYJz89ZO11
u0T/Xzu//UPMT4WIWp2l29XKcfsT9L26P2gMOaPhkesFuNRlASNQYyaYNhGqTVKHuruJyl1djFIO
lPQOVRvCcAoGUn8J0Rhiv4W/NgIQgbpHfJWPYmONHQMUdeqLLBDQyb7Yai4ygQGczJocLt30wLzr
udqVIgP3Ed7r14Wov/561CFuUd+1EtNKwWIphJAw+4h+syPKTC6VmLayMFqQoTBWygSaT7v7YI4X
nwMnFdNwWrTyTJ+WZbWBoK1HAHzkMIY3UoPY84czDZd4f0I6tYj9q8+Y/5UafhyaEtI3J6wRJzI5
p9B0J+EPI/5mQVAleeG8pZNeJ+Yh3cRtGPh1eHOFyuSXQdDKxWXOZwTpHg8LilovXt+EFMQo2vlx
y7Y6rbx4AkqJNmEMcQzS81Oeax0iAGeG3cEoqMSt/4QW6fb5L9kwzyfQU9Vzx8slz45/tRqnxg8l
DTLuhgAURJjCeJ3bbQQ7v8wLggRvS5veiZUaTeMh7soivgoDz1q++LalfElTf0s39JfIDIjhewad
IitOkVAE3ODyd5pUtd1wM8mJXYQcZMIckvsruWWbZdkawmVMzaaOuVdAaRCSc+yyr/3O5YSuH4WP
IL/F9/tVVbMSIROOATbhIOCGMLAvbgCSYACSRlyN+Nd7oX+b2drieIWneL/jvtgiUP5LQUQ6sa9O
+nyYgEbuGXhErCe20Ei2OrPSNa6JlYkHu0KAkmHg9enuNs52Stz4zUlHY/rYT8kInqKzlQYMmZug
v/dmgGskQAuiNG2MURLriiQSxRbuaqv7zPNC+cLg+WC7eVd1uh4oB7+eKmjOqsOgyqroigo4x1H5
JFNgT0ZeJ9UevOTJ3TmQ0nBdU4YYmeLxq9M9h1rhgC9ReU1eaj2NitwjwpcqUyShdGYNd22qL3gt
yiFwuVqFy4SSTT68AxGLILA6j5vkWeQGD2JEgnUwUkrnVmwBE180NukE0ffNjrKcoTZjtajokd9n
ceGcrU/kB8QoT9Ko9+ESN4lpuoFJJ4kvwMvlBxOkbGuDWBTR0sok6S9k8jubOiB4MqPjEXAyHsWp
oqsCXgITYXAxL6Pjup/kQ+BAGLNncV0Km4n1jMjrSCs+dossj6aiyGKuF+4yeUvFSflMtnj4t9Cm
Ao7MeHH3KqXxo3zeHwoKXLjCZJ8LixyRRMaMK8urJzSRA/pvbBDXE3IttAIJfjvL4HcRtrICaY9v
xwbueEP6Pcy8szhfUEm4McXoU02Va8OHCqIqEKSI+tgevIj7Rq/sIQjRZ2Pa1P1rAMbaLsxPpKTS
5HbNQs8Tkhps2RvvhwFJQDJHPgVghDylBDSCO8c/IO4INGBbvMhRdgWEdoYuluyCZyrm8516Z435
flvsvgLEYzSRcRBg2M/X3mIIXUCHcI5f1AWmRY2ovdpj0dVwZV4BVRGsAx3AaQF7cybhO7476NNT
F5qCfYMGVOhTCMSlRhQz5fz/G+9S5OGclrjE0W5peWVAwHVDe7jvVv9FwV7DJ7APYenLrHPLDUUL
ylUFG5n+R1LAQ5yR6LDD98QB5tbQFBVlRVH48s/R9fu+J/XfxXqSsuK4DrU5rQKwoRMoxlvmoWUp
sTMchUYSMn1psE7Bxq6wuYQPIVOUQSzCkxxD3xFpe1EYNAPNUSe+ai6O8AbgKTBsk9IycbqUMvbE
LqTBCG7z06CaQDokn28l5d8nYPQOD3tikf5sCMj6beNTRy1tc9XDoXz87A061nVTHZYkw4ZE7jdz
Kt1GEw3OdFxAcwSc9zhLZbs5vgY4lnflk92KsbB8tT3kQyB9vsYuGl/kvTujX2fQO9sWaALeH687
BNUz++t8GFnc4TSVxtqV8VXbtMipKIsBggchi4ncJ6TVItFff0z0xtYq16Mzfg0zgesUelIca0cI
InYN04Svv5QuB4lZ13Fl/Fv/QM7XePP4e4cLMOcrQ8MubAsJEUqFP3AZW8YXKJ4HSvjut0f5Nx3u
LwSckfQPZJri5lylfRATUgshy3mMMOP1zAbIMSvvj6/QF96TczWe/Eb4+7z0RTMFwvzXH2QkEwMc
c3wF/G8M2Xg9OP1vUdeyl98SSBBRXmlI0F95FOXr01dKY+rYCmEuygSkIli47AbRQ+4JhBEIKQyO
si8+ow+Mc9H5SiS8kWHsizvfRyzOIk+VJr/wwivPeaKJWJVrL27RzS7JcMqMcl7WEOf5vIlo8iXk
mGlF5iK/9w5guFQxA824mrWMrudnk84g9RoGwdhGw2VuQMVSGQLw/1FwPq5cb7B0g3iLa2aJ5Zmf
wlfYd4fAgBl/cTZvqRPJuIUVW8GIkbF70RLihEmWuKaw3tGqyfu7JYV5Ybce90mhcMMshqQmroVS
tX81/hox+HO2xJZ4AVHEmYMEbrMF1c4BHVb+a+kV4M5PeDiGKOer16T4CNbCGVQpuBXwm/XqtI2C
yDM4MIe89VJRmUbaGND2bckHmMObCoXXXDiqwkdX9poeCQVAgmQ+S5QZmteLLCrL6LQL1uJnm7Dt
wchgjV78nkFtlYN/Y0oeGrhjB/ik6W16zPjChSTIqzSYQ6pJdwWKNIKU8zoxU9JVgYG47PI8hgW6
SO6dsljYlDmhsWXphi7EkV/ph4H59aoMPu5xNjBrovNpzwM1efF0aak08oc+OVer9Yh66ordd4CS
GqPzyMzxGatJIf7XXvl8geWN8YKnQmZn20Hn30CFG+8nMJG92lzQitv4CwXG2qvzqxW3kbesWpOk
e8CsbbsxERFHqdxxp53ZDo4jhmzI1qn7Jhmh7sN7t4EaLNkBu/KgIETAICXpurx3vgQB954sOqVu
5yo8tqo6ElsOqi3p/m3rTtxxW1lPXQe8dyiO0MAecHlMJtmT1nFqbLfOwSJGQl4cYPnvkeGxNhKh
Q+LoK3k/mbDXpnfrRFoC1JXvMJoR8Z2BXVNkaz3Km/0HOK43q0+yCQoFJ2WZqXWb2z/gFdjhlN+G
Rm7My3zgdGreQ5f76DAGZskYMAbbCn3C6+84GZ8eF7fU50iuVUzTQ4O3UjoarZWHn12+ZlaLzuyV
AkNDSFEqd3MgEU4zyV3uTZQ5S6gIP2HD+ldGutjrPphKwXAJYtkzGzmqkMYywwSbGQw5luruGJOJ
DR14GsiX0zpsI3uELe33fRikmVTFVhutT1ICM6sQNd9vZWRVyqCADW/mo5PZnHBRHGiKAwrkZjPZ
SrA5NYJYx+ckWP0mRAnBl9YYjXsKjCHN/oIySlgC76nkKiumIn6iiJLpNpNZZE3PM6O97eWkYQ2V
OlrdTbjpJ4PUaD/dgOfxw7V80raB51+ERL6yGB7IYz5CE8LjAeyvdB/Uta6QYiqTm6RLB1SKKcQY
r0fawtiKqLr11U8Mp0IZihp5iWOPl33Ez+MnSfAQ4VQnLz1qujwUIbSfVSaGHJVjhCbMiXvap/Wt
bHBmp31Gh1Rr7bALd/toV8MHUoonjxgXo/MgOpeHQVW/szt5pwaividdiGADi/1dpAPGqdxav41j
epHxMe1iWG73QW4QVWANjbSo9X8ItE42j/cvmag8Z8y7/UEO3sZ2Xdq2DoDy0JmDmyUUclDBv+uM
4a0aCP6sYdUelTLJpuYaty+I1sZ3wELqKNScjtB6eEgibFdewzOH0SyHhBxwfsBWyPS8Lj36mL90
4iP1o+dKdVPbkia5ir7D54wXwhetMHogLkgTl31qy4/m5QVn4AfRXWPPI3wHec+HfC3z8ZUwPRir
vlGid/tWfAtCTp/B6Vwb8NAUEhnxawqH/aaobpZaSJng6PTeTMIBHnGKcVTBhjFnmiHs8mJcT/wM
H7fOAZQEqqbz4q2bKSXZ7tP5LRntSY3OisxsJIa9TBkdja30bz0uMQcXmC6uHnvEySmEjCPVnhGD
l9LcF0mMwHNRgHRnXxH1kx/+BJP3Rme6nv0/JVoL/rX7Z0f9FFIfV2hi2ECdvtY/Bbr+HEeggF1Y
nsEdENwNQVN6XqS3buxW93Wh8+tFl5t7QfpXlgkaTyGcTFNjbtJqh2MUFgYozR49hM7FIXeRieDj
mA7rZx6kqJ2Y2aGq0Li/97Td7J4DqcZMFmm5VzKnw7P8hxw0lYDQqAw12mhqhPqfuErmiccjBbVt
v6z6NgbyFFMa+17WHC5G8BKMwE1kXQw5SWOrDvnyPWvOKGldY0XRqCF7MAH2D0JX6m35/prFfx6O
rqpS5ceacl/PhWnKtz7c1K+R49LJZ+TpkBaKob4E4X3witEp8WUVKHnLCjJU68Wet+KPRYbBH8ps
TW/YYSGwUU7mqsRxNxVl/wiJ4KhLjrUNpAe/H32n0TozdPmKRAtUGqBTy+D7q8fwVTDZ0Gjnqdk6
n48x6oX7hwJGHseLmpCuPAZlfDmavR1KFyMEMEw7kCiUB4f3gJBhLeIQHmxnbo5Qp832l9Lh9Fr2
GPb9Mqt8q26Ls8k4i1ineQtYFtgleXWR84lmKKGggGKpGo/AjCISvdlf9YWT7SszpW2txbIUWoHX
bw5doKTxgUG2WrpIa8OqvwEs2A8gIX9KfkIAAJJz24FeQrfAsLZLlmPG3X3rVMvM68/0Sk4yOT4o
6QQlYASuzb47TQESys+ek5LANY3Z9huENW/LUkPqBpFdwDOJx3ODT0aosSNyYbpArppkgvPcs9gl
ApBsw5AMoXsHpv6TFMGA3g2D0aoaoZK67Naffy807HSR6Y3PquIGocFRI6Z2DwoDF1/wJuMe8ZKO
wYxoXXtOVrFPZQ8L1qfhAYkN9hLXMpxFlYn1jIYvsmPybivXIbSvRTAi55K0lG4KTlrDJoHSWqPr
FPalWoFBE7MATgjSsZBUav7u3A1asmRHjVovUvlF9XD4wYLUOtawM+momEopQIyy9ywJFPeuDje1
wTk8VEia7QksCYjiv32lgKbHLf4/7Uf/PVa56GCAL12SJnTUh/xPKXJvVLEOKsD23A8cOf06XR3q
eR5R/LoFMZ4Pw4tYBIVz+r2mrhahskt+HP42DhjqS22rJ/YFaDcngr2muHAK03HPBKPvXDfd7Nno
F8dX1IZW5thDQ8HphTZvW+D2g9816rtJLn26gAmwCZTOuGbISvXpL+gmYlu/OQr9A/+/6KCqDe60
N6XJ6x8mqrLJOmuLLHg+RFfixKWVpr+NMXU3IoqK1TeRtcgadhAp798ttR2uZIFz/XgioVuAhFIN
XMZi3lZ8u6El1vprjLqOgDQteHRqm6Q6A2PhbrGHatEZUgAIEfUZH7XpW2Bz65qIhbKa/GMZ8Mvo
Vjw/9YU1kP00Aujt3lwL8iWSFFcoTUkdxz6Jhrn0AmjtIoGl38jlfyRL4lFjObYjZY/Z13aIUfJ8
qbDoo6Ii2lF7Q20OcRkyqSNEdRzf7yXdwtOPyXKtfMqYreDeTns2MWSx94nELKlyMlJlPdcKLycE
KF7EthCZLWqbpM/mXdIEUzTMT8mn81cHzShV+3LzyEK2m7iyctKkzQPJyRACvwaa9yUqlxoEUq5E
/ZKsNOXU+4mvPWjrYtApZzSUuEuBxzvr2sL5JlU4Jjdc72wRKdegY976jewDqRsQqF7Gn2kPLZ5j
Lwz6IitrF5gztazzF/2KF1los84+UpFGFxlo2tyWyLXSWDylXU5zoy/bsH1DKq0GFIdc0J3BJo5S
irsLEiGjLJIY0n2CXJPA71EHiot4zxXO4Pwm9ewsfF2V0NtMvVemxQiAOneAAMmiWpcBtaJ1BrKO
irbq6dxnVFTDofqBLMKdYSEdKPeejVnKC6NFI1Uj07juTSkCNUwHEP29Bm8ZXq12C2vJxpaeVmbH
EChOzzEyVSbS5bSwKLaIRql11njdXcfY+vxL5xOZBJuCmrLexN7sgpVuiNfqLLAfgGyTng+LTkls
ZIw+Lhq2tRGjX96i8S6QUbfzMUg1hXpfo5cjB2y8D1mYxhUk21RU6WMc2VhDKCp4uKkDvXuMGkn4
QXSOcr6zKpYOx5F0Zqobe5Bc0mQRxQjHW1nfLH8lQ+TAWNdnZ/pcHf3hfRsvKy4Xg+WjcF7DTeBI
azHEDBM0UO3cb/zzfeQq8T0b8J4LXye82AoI+d4GTLGs1ze+gRd9UX4/IaIsj9K7b1/InOTzBxpn
5I9NBH+Zb9VIto/KDldsE00nGC/8JBLEU0J4LNOYPQPWwISynq0PXDZxyolU2VEOG18l0EqCmWGB
Mg0FcyR4e521hGjevWqobiCE1TqzKrSFhH2OrpjT2ZJXWdPoofGpWWqKQlvaKP+GZySHSZRWNQxa
VjURFXeR7iz4FpvpVPLNcJmdnnzsTB1vIbsn66vqerxWbV5XemQoXBywicqVULP4vtaeRdsu8fed
lzig7KvKpnftq00Ul3F8h+0yKyh5v8iZkRmPTiC1N96bUe437epW3eGcyBfFICda1iMYAjAtblMI
hFYlRZRNkav014qWJCiHy4jKlB/g7jd00m/6C4rZXoEhVJbeJwhFd2iXfavC0/db3sZE1fDyRS8A
Ivt8pRsDzUOBE7FYeaHBb6i+kkR/PWd4z3rAhGROGhhoYVVSoubvxLiwo5CLkhF9UrzRVb9t7iln
gGwcelwNAaSb2Af+DidvmmBWr+yW3hXpVjsoZZ7KIZCzjfOcX5C14X7l1Hcz/CEkWjfA8yg+CR9h
LhpN0WbIgeezeVFOqiqhZrlOKc7njGHA91ct7DSTt8N1ajNqUUpCZdqN4z7A8WiDfl/ze1HeS1No
JOTdxQ6/Qte+VasfNHwYTwpow5Ee9+VshXV/n8UlrSw6w9iOLcQOMyueTNdtkRguwpjGl0sZm1sh
z+zNrnudYN4d7wPLhKo4zMlHdJzygnVsOhvCkiGJ5JpV78aI6FX8LulHkxp38G8KE67xqi0piIv6
gVjKyIu/r8XeitVpIu5Sr5UhMjvXHo571luMuduevjN74yyl10hmttwOHPqE/Qkw5T6KhkAZu5sP
6hQ3QT6XNBOTokfUwfDTCEEsbVMFXkw/bzo3pd3TcIF1iQn+n9L64uEVaFekVr1djG8Pk1mVJNmZ
/K4QxavDHmHmpWpqaSybnheYcJknJHmxXgH45Nq50com1bWqHO1CMgFJAGAOcXmGncpHki8kh1Gv
BVHAOKrAa61hv8o7AJyUhEe8Lmms6YSPl2SM+CNWhow7Bc2gPZWIOK86tj5nG8MMrzvocMbooHCL
SiDxXVuvbPqhU/LduzBguD3zDzlXpli86XcJBtRrcJoyLrWxOh60Toiaea/u9/DdmcGLsHSGEtQp
MS11xm5CEmszeV43lzN5ttKGJCuWRSp/wwww7AvnKC0ch3uewNgm/ZyjzCWgT8FX8xIB4XL3rEIR
NIuJEMWfRE/AJsms0U/CVQZg1tZ1Lvy1lAX74l0AyusbtlJbkbEeafB2DX1hRPr/u28Wo1mfZwZA
7RGx2eNiyYEAnwJvAp1Wm/rEaJbM08vyS/SjclAKftkDa0L5MAEwSSVJmGJcdc15Jd24WnGjf1iy
+02ZUETcLa2YN4u3HQLVxMogkmtEfvtkmVEN/B0kQa3kaRH5VSe/z25crlIoLrxvuHJHEYxBK1so
ugx+XSypsy53KbvvTIsZbtludnwkqeMk4CNOdgPVrjcqc7bh9qOfyQllwh8/8wBHmJ9vqBngwyLL
o2QkXsK6nu+IWGj110+6F99pBxLPHLEzRmalkLJpYIQN4aq6cYSaQrcaO+mQlrATcSssJLvzkvWj
LqkBhcfSecQcekvJdQNZ0Y0FsCoX0pMmElKRQU+xCCNm149Y9lQ9Ai7bkbDtxonQKOY2hwu3pEuC
PgqzcYxFxpWkjFhm3yum24/HZ18aqLDDsa+BWWhViTKCpEOOV6Z1CCMnJ1BB4uKZvpWl1T/6W64N
WSQIQLee81JjydrL14heIOZKbEhhpYu8E0fWuf+3kydM9kaACrL8k9ktzC55bDMo+8yHdquqDglL
+Qp2LCuNtnXiuD8ojt2tTRJ/W3Wt39UY6PkuD123Mei0BUKwpzVkPzMqo66UpbvNVEwYcS+9GU3i
iMPRE3Y9h6A35PNAwVFrYSH8W+WYzZYg1Dvh6uGaqQfR2ywQ0UilbVo2KcTbUZKAjt8MGnxAlvjm
MuH1dt9bAZoD0QHJ3STCcKOtuYv24GiKHwjB0bwdOU4nHzYNMpCCa3x5pnluOQSXpwDtmvHGofv7
D288bbmJV64jgXMlIYV3D1bZmljH2KvfMcMC+9badx7q5BgAAY1qI7TCJhKRoMa6+qb/v5cvPPWg
pvQ/4i3fUeaFxcCKNC01XI+SqOdzuV+wYBwrO1uq1JhxJOwMsr6oTliXw5KowhyIJnT03s51FbvT
xJXLsCQAes2jKX9A2Zy9q43rAbCaXNjbZJNykRJd6d1frUapol27wtufI4QVm7Qud1AVO0afecQA
Hdtw6xZPh5Rbuxnw5vW0JHbxYN1POoZz3XPxI31ODYTmCIS+HR20n4wuqS4EJkjWgF1zVmNbM8in
HzMTV1++92Obha65aG3jOhGIQrJ1tI05/VPBH/mrGxNzEhK4KYfJZzEUKh6JHTat7712Wk6hQMFL
5AFam4vrWS5DOFeark32uD534f7iMPbMnOcUpCfxPQjtNOwhri/g4choFh0RAjHRkaBv1PlEbNZ/
w9qWZc2N2ERP+t6Y/izHJBS7okEcqywgBnUmRmMAFBfr1SBXkLwhQNI1iUHR+yFtCD3KMQB/CBJ9
1DfTVi8buX3XReKFymCPAeaijM8Bt79jcOdwxOxfLVCFKRB6n1yi/Vjq4n3BZ8KPqOU3YxjPicyl
me3zAgxi6I6Q8z4Q1UysIAXMlgHHVyY2AAzgpGQ3xMWboUhA2ADTpmjUhPtErA9LhFsxLuYokKzP
RGAlwhgbGpT4x6hxafJVfZzd1MWm1QIWLlqcc00eZQtnuhKgNYzC2BMsZVPXw8vuHb9BvHnyJFFI
kKrjKs4wLLu4Z40552nyzq1wbMGfZBaDkBcAV47ctB69W60BoQctkaEfqasxj8DFJPR/mufj3HX7
scissMAWKQ9+pvE1Si6XMpBRCAgH40DqOFLA1J9WJXy4xhuBpWtpsK4FsIspDckvTFFF9zjOuXO/
4Ji86B6r9yETnQab1AcfuZ3Iu0gZjMti9wr1MbAMwNixGU3k9SkyP6BOYD1T9B11B4efUxqthwm7
6JaEJ/GdjoqnGxHf+aoZWjVzNo77yR9mQ8t2I+jVOB1QILygQYCfju/sHS0tbBWfDEBg6w4t060p
ywdrXJz1zwhzJ5OTr1Ahx3en6dIWnW2HnizKQE6kR8zVNgEMeKlsf2nJIqJqSHNkENLnRsli8YeJ
5f6ka2uJYeRwh1kOBmETXKD6sUVd/XeN/1OzCGMY8c+YcBICQly3qYWwOiB+GHbrxBuJ2pQosmr2
DtoPnPZgPuAdq99QL3teur4ClwQ55ZsITUyMP+D9ggn0rLMGI0iHtiYlFwp6yMr6lCGIzM/MAj0A
3MKAgyPKdmllImOx3zzQLF55Ap9smjRTms2iD3zIdJSENM6CB+709BB0vSZT/XYYCZEIMJ4i9RqQ
V7/3XI7g+uIBC+WdDuD1mfkG8g8JCsdssZIPlj0hOHR4pk+fOJpsEi1CUraSUDpvJMxFGBx0f70w
q/7XFFd5yGw64vB5nNT3XwRhA0XZDuM54Sj0SRaV8BIpx9/tAIFkaVtLoqRvRqsnh29F/bEEUbhO
RZoq6vk12wJPaGGAlPfVq0MDCN1SrV+/wEkIemHbVNqpBqXg2S0N0EtpIunJR4Kw/5aVeqFJXZuv
EagbhBvMVjPehOm8xe0ZmHgbL/ReB+aRs/O4C3rvbCX5fP3uIcElHLdyfOxPdV4lyV1rKtkOPEhc
27U4lMbyY/B1l6YeWfH6QaJjHzkCC5dVXWXKU7g6McyKTzHa54UAI42OIcV4ZAMa4xM5q3/z1qPb
W0qp3o62tcainMYLNTZsNr2ojEQk9ruZDEvyFKGIGZ0KTbhq/02gHwykNfs5kFu5V4EZ95H+dsxn
sM6fJYjWqp4V75NkOq4Cz1ENFsuloQ7UCsPq/oL8AhxGYFSi5ohAXy9jPJtP6bL6JO4TT+S2bs1S
b/IkleNF9i6ffq+5to9hcc9h2RMrnOPFn3epqBdABhNnk+Y4pah3B6LqmW4CzLjsL67LlD2txW7p
9tAju2SqkbZ68uahBaC8m9cgTV8CpnyQQKOHTYG0QHJkmF2H/Q9ba8q5xXUT2LQJi8zyBv8D5WGf
xnzXwp9VI5MsxFRKwN+VbsL3T9D9rqU4VmsfPiQuqq6HFBzRghjzari9Zi6FeoVCUY4M5xitdzHZ
MDOxQpPgJNYgvjKCxKpCr6WckrzD6BBppIDsgFs2cZjBsKNa4tX3F25JJR1eykoEuceafuN2gFrM
GZetk9Rw5fI3XoKc7ZbqGcNRne1D4kq1kPNASvyfd2l8tH2hcjtVHgCAkclASE0zKn8VcDL00+bF
nB9BvrSxjNEP1iX9sZAVK5Ounjph1nWbkVzXZj8NgZSoa0qIS9czp2ucN/z6CWGSOidZhdQSnLhq
bup3le52WZtbB6bMVLZwcLEKNRiZt2Li/CNMUM6oLDdF4TxLLNqWtUjAYukgM3iiEkKUirW5pNJz
YfR7RWB2kI7GCWIweK6pwzeDJJ2b4Xkz3bKmQNpe6ZQwN1FSY4p8ufTt53Vg86mbxRJI4GnDLbKd
YoUphizfZkwgUCZoLVh9WAtOCWMcj5EScGM9kYhYFnXeMleY8cloxF/9XBx1d8IeKJWB5H93BH7f
XS8NKnNYu3pH3XqeJd6VOsMDNtQ6zYWMbqxRgQSTCm0DLgkqBaAh579qrytnBsJBjkVwtik/emo8
LrKCnbCf5vb6VWzIj8m8jvBT8LUqid4EOtB+faflCKherkKATQa9GpDeyJVzg3rEGohdA9tr1C6x
vzsGshMiLtXl673jc95vdw46nzi7GMieuQWTBpsfg+ZkTm/rRiS7eJJnkRPqJV7blq3etNKsuxfx
qAOS7iiUYDumbJ2Dmq3638ecEr+ZfxJvFnoEj4yqPLEY30oSK6vjy+COrlfItbeZoRxHCZFU5U2L
Dsep0YGorRh2wV6KCkLm9yqSD122ITS7UrhHWI0Uc9SAnPqNZhfpzpgHb6wyT72xK5M6dh6p3zWE
Cx+lKPrDdeLNk8vsgou2u3hHDnS13tLCtjlU8Z6btI3HQpblhCtGZSe/jrOy3yoBPkuH16wARUhY
O0KyIaAaejDaWKoOt5GbS+A61sJB9YKdDcy9hr30FnphUEAprD9EHWycTV21jXQb4cIaZz/jWY1W
NxPqfuFe3/27kGEw1Ruvxo/0WFzKZXyR2/8mWwtO5RR0/ZAYXiAp4FJnfkATVUz1PENESlLdVemz
0OlOFX1Lt1/2HozbhlpcuwpYfiYAfi3JT1quZXbvopscV15cphw69ZhtxB3MF2fl0topq/WajhgV
/HhrRvQm4vUU5IL70DRZQoyQ4RINw4dwu4edGIbBDY4NeIfoeKOsXwknEUKsGb9LpCzyGkY1VvT9
9IecwZBWEyRGKpBoCXdkSvZKKn4q0hIylMt3B61ggconBFnIk+ovD+zHLqoBJENxW8cFT03EzqEV
HS4CYBs5/nRrVQbwDcpig0c1y6IrsQDPW6LnoJWFktI7fUT+UPvlS5pOOLsYA1pMiM5rNCcIW/12
0bSifbn2mP9qPZrqD1zkr9ma/4lnzF7q0GpUkyu7Rg8hxs61z789aK5oGRgYx5YO/LEuBE0xHYmN
AafHUeovogmpmS0VYHpjj/UvT1V93E85Rp6m9AJ1vy1Xkt0XpnL/Pt7KLAoiIBGm4E7R+E4poa16
hBZBFVAd62IPbAf6ZkdWhuAuA7UZ8oauiVkr9MwDKam8vMNi4FnTFnbpA5C7+hO/kqUPt94s+jPB
SM8/uZt8DTE6qqizIhKrMsbWvAGkjMd+1KuHQdk6HIhnjOr8SM0KFcuAkUsmFBGEC0gJBAybhcyv
2R4Ltw72Jsc7yLD9H3tZOdFZpL2XCOINyYWHeJ9ayfIQ5WSueVfSBGk7L+22Eok0N/6XGoIa/e/D
53PGAIcQPks4KeKY57QPKnCkHgqZvSZmC4vgELW117IrTEMr3tGxiKcJhiHmjtZpEv0SHN/8liCU
tt0ZtmHWc7Pd+AeHzqpZRaS9ZnVauDbI6upXHo3ieKO7wSZlN0HAzCIHOkShaJYOtWD+HNVgTcJR
P5VN0V7mku8R+H2Iz1y6jXk5jn3umfG+uakGqR9vSWtJOtwFw0ayRpRMhm3FhOVws0ys8CEqDdHY
3BnGFayUkzCJHVis5JIYz1NtsC4s/KsV/lifiIRaKehirzcWiavF42zRYIlhNJ+ciQT0m8l98dGB
AFVlgH5I6ljJo10nZKNpDPF07QPFV2oGmGQuVUiFj6xjUSHoe4ddRZ4KDki8C0lMer2OGzn0/mPf
9AKt2axUHxWhVf4o/H/SBdDERqMHlTlGJUYlGilyz5dP6Wkaww3CtLc6xmcfJtChc/ZsUlnQNtZ/
zb/aIsX2CqOKB4GJykXsFFYsup/fpXEh3VFjsuJNYU9EudPNWfC1EkHvkMbiF+lSKojP86Am/x+B
gx86Fne2edz94hCfyPsowqEaMMitXPRP9JdEL4J0X3JU+dlkZyNl+hNI5BSwhEPoZ3lyJhL1j3ph
qImJ0ZmCsV/oFoOGx8zZCBVfvip3ss6D5hybjvYtY7S5MkvTxH3hY0oJmsSTdvuzHK9RsVNFUrnR
Tt6xKDqwJf5wN+2jOhrgX/z63jho3S1uDt1jj43oujqwOlw/2kdMINc4/xYkkLs7vQfgeWQj2LAs
nTcBSGSpBpq2mESM/nIpO6qSWnheITFYdYf5cyCASLpuD/gSjM03isqk1v1NJIMFZ0TQlZQgE03M
tHzEUdADB+Qa2p2PyXozdwX6r+01uKdNgc5nvKpXpiFaVtqcVXyIFOHaGP73a8uj79y1bRxpYPsg
oPNaLVXNeukAzm/B+rskU58HumeY8ClNg08JW5aPe1TiKdo6nu+UwkNC9GX6B8CTXRMcv5Ssjhz4
rIiaMWiuTit+gKPEePaFR00ZD7kV3PgOgn7u7hy8miWQwhzT7y3vdLmqsk0lzmm11XojrPaaIszw
qkbBBmiFFILqb1nh+Ntp6sYmsztRvkTnuNyfoboFOGO9GQYa2BveKUEIbOQEbxLq1WubWO4Jmcb2
FM31W7sjgWlJGmhGzehvt8WeaMpv1uSO2kWomSjNvLRczp1DqNIVJ9dw8gesHgXtSXXtXGD/1QP9
WIOuJOm0xbLfp3fCurBhnrc+RFolv2yrRpdhAkinx5KpRKJJ24ffgHRqegKC3d7uIi11GT6H6FjC
sgjoQKcXcypsaVNmbokTKwLoFVICnylGeG16IvPKCia1LBFqgj1/JQccaAKH+xeMhdFU18Uz6hgq
Wl0N6x/EgTOmeYimQJw2HeN+GYjOIjcaxmjjEC/QmB/duZa6LmyWjyyx+Sp6HpARoM9/5FO6JfMj
RQCoLGITklO5Kza8d4awwqrNwEqOnEmrJ0p8geJ7V6CbhNmvlyyR8k9mAGJJFIU3KC1b+icQPKdk
7ghHPrNfNlsDTOV40H5JBq3bqNG1MP0/K3BdkXoptJqr80ZcslLlbNc2Mh35alxbXVPTvWuTaVDC
5dSGK62jsHCkm8znhBUeVc2UTXeqZmOrAt6TmiNCqeH9NVKpO8hvd55ZUm2rTQ6Ui1Awo//UaVPG
Rwy0BvPxny7wFWnYaocBYqDJt/qbvoG2Q6upcXSbOP3pvhYD6YuD+p4pbBxuKhx9N2ZQqWWCoDGa
7yGbqSWvyixtBfovOlCMx9AbTDpHvD+xbE+SHrd5srG8o1/Z1YRi1YDiFXECVdFP3XmE+9VBMMIR
gwfHttkwPEo4Z2k9Scy1Tzicg/Ne39d/GIuyJQaxjrOCq/sTpuyO0Wc5wB3i6o7hMHt7361DYZ5c
69Lwwu3aBO4VROLM6IOj/TkoqJMVN2e73P4r3OnJS2xfkzAhvCqt78S+brejSqFQLmI2t1XKkpwF
4uLTuWnhX+zCi9TYI7/j6Whad1hqmV/na5j/XQLZudtrg1ROds+hRQ/gK5TaqlG7olw+rnfDeuCI
XrxznWV+5Ej/7AmdALzi9Rsi41xFdsqnw0yh67KyBkHaSdgo6iIRfewSL1oHFN33OWJ19/0YsrOw
lvSdFjk4DW7nkuB2KdApjii8uz14LTBQpXWFT2uH19s6cSm9GD1FlvIoGA5gXSNWsyviAWas2wII
gZUd8W+a1J7S13Eo7CNf+XhHZbt0pThT24t8+uHeKSKl3Q29VR3q2H7PTkQDuXwGs9iEs3FCjAMs
PSqC7tFWbmrBRg5f/0Eenc/uLy+Lh45SzGAVweDdov7PE80YtLe0SN5SLS2SY/yhAVz4fmtARdK2
TX0vtc6lp5dF6a++FaCLbzBLNZoqosDH4mz0KwrpQQ7+pO32IcI1LPXpZpKnHk9Ag++Wsb8WYF9X
+3LdrVHxQoLhGxeT69+EbStQQfSKqhwlBSNmmZDovXeL4Paa0T+iHSLb/PKzE5jkvUXFiAcXXlwP
Dd6teU1QiyIB9jdjBj2QxMTiSIPfaUdXAwbSCilIoVt2DUsuSANTcnKHEFMBNJGzErR1oxzGMxil
NO48n+U6DEO27VUvEBago58OCjxcVtKq7SSQigk18LqRX7CAQlK/xUDfjxAWsBMGwU4ytLewxAbS
U2qA4YCFeyyi+c3SzTUxc01uAbg7aajHNxqPxiECcayqSlEEZKQcafXicku1Dz5yj0zgT4j+d8/I
T6WX1/a2llgz6PmaQHyLQQcKnQqjh0a0e1OncXcmThNxSU/rXugjVlJfHhha00qKX0CCj4aAGFaL
Q3nxsxn1G7E3m2WBeTAVX0+I6AigCV5jllXCxWeggh4W9sO88Zrlc7YWwRVf6iV1d/Uu2OVZydI9
aF3QEYKS0UnyLjaeHxLt2M2cvtaVIyZBAMz0f8rqPq769V4LPYufwo/zSUjXObiKxNGWpy7b4dsg
s2s7lCXHYjX+EqFCN0HEGDdvR5pUhG5zI2Y0YAQt6wKcH672J9K8Ymnqs2y4KaC8/w0DfFr8A602
/00s0hiKlqQBv5fC3GoWQeeYM9uxb70Zz5SHZVQ9ZYR4tght3zK1vUUtVyOuAjYTG1gemv6T0aqZ
FhGo3b/9MEoYGmjubTaUh6t8sgk54dERm4JyaE8/MeQ50bSdGJg2Xp1Kg3eJxzqr64h+Sr3ekpbp
9SUjhGPu3oHAmlVlyfc/IArNZbCW0qgoXAsRDZrCh+B2h/ml53AiNGTFyorrqrCfbT7plaoPtPq4
fis8G1jepuf3TIHxJjrFgjHv2ALVygy7EIp8yQZ6IP118ogocwpXivIrZI9GK9op7ju/rE9GSHAE
SlUZy7QJ2sEXNlvo50t5X3poO25ZU1THw1C4xc8tcmGLMRzYJFQvFfZ8BWuMMkaL0KVC7JGmG/5h
5FDO3J7e2gJC9kApMTQ3csahejUocXWKGsY4wIG65DSxiztpPd8lZWuxFvasCI4ql8MxTEguEr2Q
7hyqtAJdjvPoMcITRgmJ3f5lY4zRXFAb2wf+iPewAs8TBynq8BbaaBRTi1YFcQyVB2D7LGgPAJYx
Dgh2iBURtZTCC/HixTQqlnCFKqokrVSw/u9vQ6xolPNfvAwWeHGer+REqltUllnSWftJDQR4ud9D
2d8mKp5GD86cWPh6yFChVhsEN6Xmg8W3kDtWn5fXzp1IpUepzXMMvsgGIJnpDidK+YB+R1941PEh
IhkBdnGRsNORo8hKXIXo3Bk6c9IQkOAdZ9CubHYwym+LSHuJIL+YTF2ucB9S04uejiDIdY/EkDFx
gqz+c4jJQK0VD3zpol82e2bhOgWlOh+GZhUd/20K2k6AmiyyuZafZ2QuHAA8pVRmk2jZWrvywR/+
N59H6JA6/5xi6AZE+RCFY8uofSM0wdC4vPdO2OgBU4v2eHVLwqPjazRbyAmgI8YrEvd4P4SIOimd
xONhHsjigk6o2HiceCNtaoWtoIjeJvxhkrcKH2SHbeObeWEymXMISgzUn0RzG93kAfnx3lW1mp++
xUbztMVdjvKCo626HH0tQ6rqAVanwQNafTCHBrehrOWxNrLazTMn1pWhkb582CIv8Okqe7FxiYSV
Acuw6Nj6Tw9Ai2QdM66XvO5uHS+09R7ijLdhC+1FNQ4Av61cWnX37KDDrx6QJJaUEKbSj/lfgb8O
WeWSyXFN+no1FZ+aC3PVID3wTiFDmt20S5tyc6zV8XmFcT0nwJqMmrn+3J8l3Tb8/b8YJjdAM8yn
4tNGG9Bm+puzMO6gJqdJBmYeYgBi5MJtmcLDnGvqWdNXHxN2BBzOaebHarww2kup26OR7aTdYeRn
JkZ0E6DuWbCigyuwYa1c0WoD6/yAH9QTR4eGx2m/JBXKyZZAvYI7Kaak3QFe3bBresVHZuL9dru1
J0EuxPoKdorRxfU9IskZWG8qmlLt1aPErYFqRSkAVlz7AvtEXMZFKbKNiDHqnxUzqwCKgYw+ERjt
P3zWDAK7zoq56nJtx7laBpliHrjplWL0YzK4XuklrS/k6M9alZZzPKl09L3oAIw8RQmnyJr1EGpu
s3KZwz0oQQHL3LxK62hJDkYJ68eD0P5xDTqe8bQFAo9o0xQTDAzm6n8EOOdyXzJKXCWHGEtAyZfr
mjSEYx74336vE34bikjW+zBi8JMHpJHAqQ5B9CCAZ0h9QlOrLCMc51wIqro7MQXGaIfYNV3K6kAV
ZerQxLNOElqt8+rWkI6EuL/27LR4jVU9ACU9ohpQx8lCOlKyF8FzHTDPVZAcnt8y8qXbU1IumIWY
zKj8nYq9nd1HuiMytmLrCIWME6YcLgDhabChs56v4zPob3G8fTTUhYiowG97ZQmMnR7qycr+sj4v
3ZdHqbq/H5mUKILHA2K118dYp/5+ZBmgAFsgWjAsS6Zc3gu5euKxtivDq2B5PTNjlhpaLTVrGSAm
xiW4RQ22uk5IfP1mR7e9OYoggJk3swGJn/BecbHusp4G4R82rajxkfegPhm2Wgodnr7tiNcWJAJ9
s1RnUsGNkxrag1SXHoFv8+iyVBzIsfn3gLId685iDfsLIoj7Le0booT51O/LhdT0AMfAQuKAH50Q
Ep7pECK8zO/Ak9t7cmEdZfaMh9rLFELBeBuKD7scnXpHqrxeKVhn3a+u561QksLbr93iChCFwWZo
9pjP2vR4nd5VbCJ6X9EChUxcUBSn/vYYM8282+/zmOSOalhnHhjgnOOwuSVkXBQmmTPlrlRDsDL5
J1LIG+f9dnSMCW+bKawSJgJ1YfxFzO0QW8ZPAvytPhxWljUuI3Ky8LIsBP0ZLATcxnDJDQhc1nUF
iTqghd8WxudUaz5oyEEELPJ5CQycUHceyYsxlgSMTG9eR6MPQcDnOR5h0cOXch2+FtIsP10lwSw9
j1Z7ISkYzG33qrKEoLmk3eNNKFCecZRZR0fibyrzAqZP4RegQZYzJ3oDS3kXfvElBKOOn5sebZ5F
PTDtWNpVPcLNewQAedLTfzar+hW426Zaj60ZZ/DD+wAouw/uDDBiv0HwDKpuwk2+j328lWp614px
tI6T4+sCmWh9XJ1cucAkCGq9/vtGjsxqB7DqKB3Lucw8+WcTIzw6Z13e2ni03IuRCYcEm1LQ3aG1
e8II9eoZJirCQ6CQLKIaNqyhFLixyT7xsLHkfKuqm+mxwgg5OTxg2ZjLYh78xQGKFVZ3GmohHCN/
i0s1b6ajupvq7zC5r45VsWfVfLJEOJxZ5w4/7cuQxps7u+hvdqlGFD2HGhJW/42tQYjTrI5tb9/C
TAG6kFU2oScS1nl0dFY/vmwa4sRkc8oRfvi3u1T7nRZOF4/jOJbkYjym2ovtaylBSjJUzoACFXoj
gPBQ1S/i+JlxxZCyvnPiuNsqFExjJNBznkJ/Luc5Rlyd+YWsWW1DwtTzylP4qvm5wH/1zNx0uENq
PvE1ggcavEpfLf7HnlqG2V2IFcCCUCcUpIwWr/9wxkanvW5fZXO9b9XjfRGzkfZp04bjFWeSxkmM
pKnwSmCOSqsWcG++3J23x88OcxRHvJiXeJilI27Apf3hQ4lqIPM9BtIKoGBX63eZ6vUrjP2QUvop
Oeqzm8gbx4iwM/C2xrmpQT2AiQXt38Tzu3rsVsxTiSbmfWjdAS2OXxfvufWumUqBewS8C3yv3TNr
5AwsHDLodHY+L17KyEnf2KbAoMKQqYUbx1QgfEVAbVTwGnrR3z6izExboweqjCvEeYuESTnCu0d1
dy5+xoV5tPq7oY/8lAVk0yEy7PvU8PQUlZ94E5MxrjX/JDAIiynQc/7n9mTFBvJNaT+ZIF5lwmvJ
8AN9wDyVmH2s3kd8QtoO3G6JKGT2FKPHdznTXPSL5++K4QMgO8DB9M6pSE0RmxAQ6a4aEWMGMUKn
htRH3q+NhcPPkw5og3Djt+TgN8qQ+0RW0Jdn68lql5+Jh+yAzKps4frc3kl7zjJJQ+gKitQfw75a
Q3W2FpPxvbceFyj2NXixkfRbka72hfF5EvrbW169ktNu/GldMirLFi7sqrqMfc4E58YSqBYII0Ih
MbXoDFsRMtcK26ReZ+mdZQxC5rjmG/EH5gzBYgOCFbpBEvcPfmF6/Rlal6D50Grl/4yKfqwRgDKL
GWDS9VtdOnl8wtk4DIeaUbf3lIHKnLbPuSRPVLuKtgQIyOiTIQd9sW+koxH9FkxLOBBmHxKJ0uWZ
lt1kXKdNHA41RZZwtZANRiMmF2zGCis3xM/5yp7eLtJdshN3/lKNSj8RPJJoWG73WJTuErVrOdXk
LqJjaao/WoaDFyZvUIil5DCflm0GkSVKFLcURL5FqhS6Ov+t61/O1nQBdJ+5pj0zDDYjFM2QVkFu
vm+gvShyAmfUxaXHyloz+KEzw/e9OrPNCXQncs10SmmbOBkpAZ+VhPNVyDhf/cC2REsGbh6qwJ9z
rON4ExI0Af8GsTSFFyv5PZfRBNVdkDVsR7JJlWUQOpL0i3DPW/Q0/+bdmdOxikEI3v/esN+EEdU2
kY+ENALqg/YvaYv6x+ChquTbfOtmObwjrzcNcVrP8bgQozc2w5pEcT1YyJrfSheokNhlAYPP3XBb
tZPGANxM/+h6pIZpRqCr7/qLucfFyYrGdF0WGPle9U1803PJN8lrLIzErUp2JgmaSp0rHHLdaq+u
eubt3vle3kcBfxUMCxXwuW9CzDsSGBEq3smgebj5rOgNXK9LAIVkYVGOCMi8TViltSXA3ds9o8TJ
7IOcujzWy4YZYAZysoyocDgK7OeqUAky8/M/w+toOQafooscdazfdHgihtu2HvhZnwAR0cL1QIG4
GZ6kHHnKAKB8vkIZ+bAu+37OUhG1KaZQruPvXYvnbYzixCPKVDBHGTzuS/BcibLMWeZNqdmPVY5j
AufgXsmqLVg4yMBXD82Dd/jFamqT+HZ3nfYQR6InqITzrFyo/X0UUrh2yCjSyJ2z+7GD5yRCcDaC
cK9S5miYvumCSyqd/2iR1+o63FPq1YRzQJpRbou31qvAJxNW684Apufqp5XRZtyq/geltnbzB+39
BxtstYGrxcRE3hmpOGBPoBUa6vSc9MlyRrMDQMgPPWz9cpYqU4Y/3CSEmuYoxAusAgZuAiUypQZ/
3DAT99Zjw4ZeeJqrBIOHoNeVl7SCg9dSCXQOGSDyLHSerUbK+JTqzSUehSB5u9wfgOFvYm5MwNZR
tLj27LJf856o4sdvYhWjO44OTuIOhUP7BrTUpnX4uS9Q5Z77jTcf6N3ok42AL5G/Bs3tIrK3/5TR
zcQMjfHDEJRfNJySMQvOv/InhmgUNBAjVMr0QmcAwzZdqdA5n23XBoyW0cM2VBLh8JhwaB0bDJzV
vhO4Zh7ftsjfYKs3PeT3iYYSzC60L+F3Dh+eTWmrHZt01VjPBnw+0QJFkMPvo9QjUW/5U2hdvJKY
4YezWdRcNT2QoBcvuFDX93NBLLOz7R36+e1ZsyFSiF7+iDiCC9hW00o9mB2/z19dWLu7AgFRCmNZ
TBOg2/33pubDXbRMpsqprO408kec6G4pa9Iq/VDYlLERUzy+sZNJJil8ohMAvng+F+HzKvn24S7r
s8lHedZ//hY1c+1iiIialOqstmZUL9UUX3gD6FoX0uTJUPTDkJSiBDOjF/JU+jtPCNWIwlYiMTja
b9zv1Sxef7MdZjg9ZLAYffUnEAwMQ5z4GQeE5qR/bhZi8iSLXpABGAln0nDeU8Ink7oUQg2NHIyo
uV1TbwNAilUGow7U9+MQzoFUdc1L5nGeBWi4PuIcV/8/4/0bgkPrllChkCnaUpuMygX7bgYOrsuq
7sHkMpCRIomNv4eCgaF515rZQOzdr1awaIJv++h3m7kfPEiBD0A9YX+FbhZOD2qUV3UL9IHBDPNV
iorkeEyrMKP7nufUHFNs8t1MF4Rui0y7W+mSS9KFdg3r4+FGK3JKdijS7QAckHh2L35bixpNIp+v
YMHT20fy5uFb9tR0uHAaddxu7qOKgMOOq5CmiDEwEF77KRHyit59KAoIekub/fvklgQOu3eG/x6M
aspO04iTgzPnBRoSMJDjlbztXkjIVy7gqrkH0QWiT0k7UkpllViRlNUndmDGgWpc2Xor5vL1KxRG
MfunaHJvEuAYljCjOve2uDGZa/Qa/y+4vhfyO2u8r7H3WN7WXaLw+z8DZ34e7pBAwcol+bcv4TMC
c7e3S+NfeOrff5EWNs1uhDElSFgHx1lJg/wIBoJlxrlI/MiF3tr1tVz92oZZR9MZTWVPE2rDDEZD
zc0AAEkQGyFVj8toXHpTqawSq5Y8CCc0zLPSFhmxn4KxWrwlMAfZElwXWqe+EQ919o9PHkcDCDNf
whc8BO6PhT4RdX2UY8qN+A1ipuX+campoadTMkyS3nQ+WiRo4ZN6FKSaGodDwGbbE+c4aSWktjv+
UEB45gD1jWr1zan1kUnb9sKLT7zrRM9FndYFLM3RgG6/v7bPCiBlRPj1Mhc/8xtlPwgCOh6lixTb
CCe3UioAialQfO8ZCxi6xqOYCcfN1Gui866TzU0zz7fBunATcLiX8geOp/GFk+91ZDtL8fyxvQGR
adNVpTcPFApTvH7qLA9ggxCZkUzSyMtPwCTTyqOM9iGs0Sg6ZGEzJ60GIESm0iBrq9iSPMc+42uM
MymZ8GWhHq78mSK6xdJPzKFStt6K9BBmi899ydIPWnWRnJnSr9RoaBz0eDXKrwkTe95RwlFlkamk
BOCWiJ0nScS377sYkwu7QNje4PoPlirlQJuiaXmeoixyzzTo982jX3whhbRtwhD6P1OUd9iNRMFh
IUJNr6emvScVF3eloOvObu5J8rCk7EFkVTDxO0BVrhqj5SwDygTsD9mvy0QuXbF0MUxSH4CmRtLD
VIbyopSJ+oguYFZH+swNzQ5ppu15AWZx2M5J9M9RWZQ5MaG6XZOTiaMwBfYDddiinx3pDJB8yg0N
b+prKkFvGL5wcWL9F4D4HvgdStgDka6XnmG8bujvjyucTp22JEeMfk/ZjGQfeA+2YUZkHgZhJ5MB
XvGT3Lb/QhlVNg7W8sBBqIpi3SS1GWoKTlDmZoxZaRATbV9W8q+jbO22wGEby13iivFSpR+SW++o
qrVAMaGqGh8JWTo6TkVmLhKxZk6//Ovk6LyzVIw7eBUG2pe6A87hqieRGqPjvDa0uKotOhYsuiaK
hBGvbPOAL/HIivd3iGvmIw8vC4HZZ1Dj9dew9ChoGZmZfj8hLjrEPjlhyUiBRL0/NMU9xXFBwgwF
RoKDd66cjiyrQUyit41uMj5/glmXdb1W3ddKAmvQ402W9eJXEzxh48OvFhSHQUce8SwVSXBCiqjR
77Zd/yHF+OyF/3kSZdPTeVr/Tmz7+ro4oGtJTyc+wOZ6SVZp+v/52lf/TORppER4eF4ea0KC+Sh4
e0Lw5Q83R2drZ7d+Fhd/yuQxPbZdZaBYi5OSLseXInb36OFHmzkcTApoOnh/nynI31Ym/E1jJnO4
L9j0aUmYXP22jn733bz654XgtmiGqbVHwOq3bK8PcH1/MkVjxupthiKLcw77RfalgSNlwROfa+Ui
ULzigPAOo2fHGPkhsIqlzm0KIFh7nrugn8BAAb4WOSEvok1fPrcGSALB0w8KsntH+rzIZ+hYzZE4
QKSIbxh8yTB/BaTCP9KdHc73SsZhOe/hY4QVTOFSKZCrKAQaNDpkx57yxSKUabiRORZgMPrXI3gs
JPxf2H01I/qZ6w1Gg9ZgUxPrrggCg4+z0GQ1DD/kCqUQYQcVeTcNw1iUGIGuz5uJRYf5SXwUOWNN
oGITXxOnAbsmx97pXrAsVZKbnsnkU8PiPoKraadJZQkmaGHtm5cZQe8+QkMScOev2+Sc/kHj7qEN
NwqDgeb3VB0Dhq87h//hamO4szktdYpRLV6rF8diXhMAdsIJVMEPUcBClxbHI5OBDL+NgDiTirpN
GKZHpc6+eoXK/aWdMBUBPGx4ov64+KjGYhIeScMQWkBzQG+97Y5XoPslql96Nk2I0DfTt08QsQJ+
jNanILYHHg/k/jPjAc4Q0PICWCsfRX1Iq8Ma2q7V9Ve6eopEc/RiufQgenz1BgFMofFZg9NAejkE
eMnrUB4pViiUZfrJQu8eXv/CqkfOMtNOZILFX+7D0D30w15ZQxGNa3QY34rsL5A6DyRfNv5wS2kR
b+0hcKrUjNF/LZYI61iTACbe3OekuyNKnCCMWQG+vMA17bzdPTP6FzBnxBFnLbTgmgS480euXSEa
t1Pgw6IgiInTgKufIp2JwH0paR39+wPzZKVUaPwqqQbArElu6BqtyC6lZsIepwrHMltbc/GdwGgb
Ho6hScx0FtElm2ALGjStt2dbUKhoTH+ylIzFWqcVfpR13TEr3lDIJXzd1GCrVsr/bSc9WupvSKm+
JmPNYISSNyPO2y0aD2nZj5gTkHR3qXDG3OrxQFqwQkU8G/n6ZuGLYEioxUJZLduz/6Fb7VCiK7vM
8DlMid8Fl+lFilcItD4KWzzo7LRZgig6yBCmaOk/9xSzLF+qAEnl6QnDfNctNmZUNYBYzt+sapbI
GfNlXhv56wZqSPPQygp74H+IKrsBbOVTpcHM2akMgheFd6BmwtRC9cFwFiFPMgODKNJ0sZMw7AV8
X2D5nFe0NaAp3850nbF31bSFmOJPrvPtSUZkTM+Wdr7mrEDLF9/kZW+qiPD3AgUNsZZnTDamfGyw
CQujUSwOIdpY8t3x5qGumwBGt/tJsTYa3gzJCjH6WpIqpvOvr6zxG9tC7z3Epxqe1AOWOhsHyTzx
7J9Yrsok2IykO5rsjE5ZeUfna1Dpz8WbezNuiLG0cOc2QvmgyeGptkgM17oSFS8BwkWr/HqZeHdw
JbVFn9gAbtTCz9hVAQ6fnZoKhG9tSe/ab1wCtIt+yGkBMu/q4ww5b5rYKbPAb/vJFZHeJHwKgGq0
J/0Zld507U5e7UCM3g+j5+7Nfr/FxdKRW4tgVDJLbXCWr7iG5oD/YkT0f08G/bJwf0U5VtjZ2+YS
r5wa2eoqa7ILqo8ihFG+ms1g1+HrPf8ZwkatN/Iw11ZZYe5xkBb8J7nWfmjP05iy3JStMWUNubvM
a+4P1qnLhWjN8n0b+n5mFg+eTuzRQNavjXeK7ffi4XT7rO7jCHy3/UnlBbXCYZnec/S0beNjAasX
4CQ0KDXpS+Kbhp4p8eNH8Nr1JzlSm7N5A93kAABFuHTRAzuKWQxqM6EstKyQl3IJHN6WrHrzpeFQ
eCRLVceOiUS1KQqk9nIsmI0QvcqAaGi+m2qrBHeyKGa7a4BDqfVuNXicRtRsk1iaAQhk6v4W/NKd
QkoA9ow+TrQHSvtIy0Hsh9LB4rpeUeeO1CLiC6wC37aemu5axvrMy+rBZUrAeohcZnP8kkFV7uj8
V+VcXXebSQ0e0LZsjXM1VaC2bkuWamwC2jXBjP5YNvfTQoSJVvLlazuWpyGbK4G7JE/52L9afmxk
ddXi1NNJjMulUDJmH+/wNzPN/zwzorXvc1eKNTsTfJ3jIpr/XCwAFxNs+Vn1DUWTNK+yRFNieUp2
dD+EZPxy3ftAlxjK1g3jZVlbd/dhOqos+tIHqU0H1fIJ3vc5GFh55dl2vvb2L6betBJMdVfucpqE
p4Q3lHG/j28C5m0jQtpOxGKsBrTq5f7RdpboaDhIf7aJOP+CqA3dxHcmcarPQ+fc/HhlrwoiEd9G
+Xnmg6EBARU/EMIF3Ezrh17aZANMpjETr1CzUmUzUnCHWPFZxxjNnGMCha7sEk3FSxB1TpcGndS5
WXnd+Yh42Qj0eiCD+aCSEqD2NRKwkGrnlINe393fiQ3gMsCHYBhG9pBPgxLQGfBjaV+MeZNSx+6b
RJxuFNofnLRx9VDgVNCM/MppaC9czpli2c8zdG6uDEnUYgoOj1BdkDjfW+F+1Ij7G87XEkSQPcB0
x7zRwC0zpdV56LcUScwFEMjEL9lFZYQQDRQAiqt0nTx1Fm8ix23q6m6GH/744fDpOoY8rBGSUlNT
F4juCnhpEqd0F0AiDTBrgdxlyO+gg33SNp5OJDnqvliDCJrAjPWYCZnn0me2dH0SP3l4tOBOjBaD
r9lCtWBkDjV2p4XpAefI5z1V+ysP59frpiAPXBlmkgRijs0b1DiNHxjA86DZ/OIDZBp7cgiI8W6S
qSeey1Jar4QxaFpPwFVgQLHWNmuIxolE+8zptd+8uzwjQjM9QX5Asha9m0qVQmO02tyNKX6YRMA8
+RP1ITzeuBhq15f91qWs1bPdOfj3m40Tq1L/5gMCrEk6xWU4CGs7zUSoBrZAXwf8LikbPLt1k1kf
amfONu3BJNX7vlYSbtqdnvoWAFaYKUCpBrB5UTlP/sKFRbCsONO3/9pbV3yjbq0U81lSWIJ2XzUA
khgLVGuMxcKLNgc2Pjt0xQyIAXEDvLsq7AGV5FkKMCwa8Pr5U+9l2cGD8UNVMsDkI65P41KFaD6d
BBxjcHQAXOpURCyrYPa1U3lDcu0biUZRZIJJ/5gVV7gqqmpTr8qgMJefXP6IN7jRI6aK4C2n7SVO
L3U+v0BvcRnNX7HQuI1PKggYWaIKUCKA+cEKcP0i2MMQIM1WMdkdI1Z81pSQI92CjLhVoMi8YVDN
mK7UGSi1olH2jWOvuMSMh08iCUCnNE7SvII4hmU3tyUTSEn24al25lnpzkOYuldjEJa+Q7TApstX
fFUguYPs+7/2t/x6r2g1Wb/stcwxivB4P2RKJTpoXOt1RBaM7gKROJ6LLKHtc5pz12+Lpgrqx7fz
utpzSnwAfLK9XzdkZRLWB1wkB5lVVs20udwcXrLSTZGRCOMoJ5x9Bo4GA4+2gSVcAVsiM46Zwviv
IZBelg71loYj3gA65vl9sGPLv0+tGQ5pgestmHu1W0eKHRRcnBLToEUv6g3LFIvIFPIr49EgBcbO
xeWFSiZ1yYC+ZinQzaS7I6UYl1Vx1KzenMQVs/+AhN8FZz7SmWqMmV/UThR1bj6doNPvP2HmLPEo
/U3IqA1lPivzm78maYE8H7a6l1HHZd2unOuNQjNEhUxnlaMzyGnnOLJ27xdBzN3ZrzDrivlhKA7u
E6RElFUlZVR+G+TWJwCeuEBHoAaXacKEjtmVY/tcMMljPVah5eFDdgPPuwxT3SxFK3d1QOdL7YCy
u7ypqPvtWTEPtEQr2vgC+gjm/g74lBvheONSK7xJsW7ekS1zt1fgfqIhw0r0Gam0jR9SF/k/bvjc
/JdQvGqTqKGwUqgQSSU+6nimYnLo4vh3IBmAGS+wEHhxaDCYEHL4SzTvWdJO8/zt/3iork01JVqp
Ef6rNdVzvmRRneG6Fkq38mpDxiQiQdhZMLhtK5hPXLbuAaDs2jjFzDP5ckDwP12lj73p1343Cib2
Oy9osrOJXg9TTYod5s1Vvv7uUuBfCrP4rc2sV1oMhDqalpYg2dIsDYLiSly50Pp8nWxFrvuECQGg
eIRSB1JtWE0GgoB2mGaIqma/SGTQTxjzZcM1iLFWRdotrHfvZnzsTJ9q1FQ5kpsJfruI0z94jzTa
Jx0je+Ph2BsmmRAyGHagou2D4JFDfY2bFpWcwAR7TP0knsLPxPXkztnwiAWyX+KOQUeZZoGD4psY
x8Yop+t5InjrSISG24gp/ZbKk2lMcHZs9hWVnmqUhG8onT6EodmBnlPkLsVKpwjcgI/waYIJN+2n
n13AEpND1/KF24P8GXD/DC3OnS8F47Sri/BH2l79LwMfxW0/Fhi58v5iagcZUk6PeqCye6Az16yJ
6gjKBAIZMDJm4LXfohh70TntXKlZzaYUZmgXfERPbbXs/XjyMtvLrwlbn9H48AJlprdGPZM5VNBk
4NtX34dKS9ln0sbct+ycBhucwthJ39F91H8BSpDwJsk70ALBb2oTeYecoQ1tiQYwS16uHWq/sfLy
2Ld4c+RVgKcSX4uA+/N71IWRDQKKnHwVHrPcSxX5pjV06KKGTCnKrmMFSbl9PAS6RpHyAZrZo8E7
jIemTdajL33sbNp1VLoo3CXwP77nGvexR5x+RqcschvkpmoDIFvpACOctqmFlZ080kpDJvpYJFLE
lcZMUR9m4FI2u3zQhkBUd+yTdIGp16ztEKPbFk+tdnFxtH4tiyND6PB20WkSkz0g2ZBlFyqbEXK+
xskuHhWSYOdDD5q94Dxp04I1t+84XL10LmtdpHqpbDB9ogLEOOvCttY3s7OyT5PFpizAReuTnAtJ
Gf9vZ6sGBaJF8q7L1uM2c0iBi9w0xmOBSsA/RxM8ZiVP9jk+XmEyHP6qIMi7vOBDsFaxW4p19KEa
4jpGqcOGJXbcZijSzCekGenK9glnvkCOw+L00g1g0H++IahTpexoJQFKPj+NXtOhf0VoVcrdGs41
OVgtLPciGMPut6Cyhz3Ye0JaUJvlkweaBCUGJOLMuIAuVXcgGMwWVjMiqUKtuEChyY96QEiYAa11
FZeK4/6njjl+MugLLy/Lil0w/TnY099OYW3k+03RUoe+VU0fVwkb4WpoTSPedYlk/lbim6Qtwopo
sM8VsYhroFt3LCmlrKRC+0DX9kKUMkDYnluM7YGY0K953pU62CYrFcO45QFHax23GsoC4R/3HYVX
o4pTyYak24D5X/+UikmxIaJjdQY9GQysvDepldFWTEJ+LIAYhmsong9RRDZiTPMZLWY9RagC/ngz
Kz8VN7mocQN7MJZWiNrQaglPpgrsjSw/PH8yunetNehIgVy/P/9SOyTyWpXFpfbjcfpB6vOuSPse
/nrCpaePRoGM2henXpY6R6+pOnfCTuwZVXGhGkNY2Twv6xhbadJU8zC/XLq9h67UJ4OVNkNVKVQi
eKpFVkvgKC7+un96xIsnrB2tvhX6LTirX8M/lUrQ3vxm+CuWqDU4mCwRaotL5E6/qD9y4bRnwbjq
sQ81xWI4sRmbb2jtWgLaLcau8Zp+B4p35h6SpyOvnhQCzYSzPqttYdySz7KpG5dnpGKlMPE2oonT
sxOGgoJ/41iTfXoDq1KGVQCjvCJYMRvLKkA15PqMwMw3bLYsRVpaL1lpW0Fd5pfB11ffmrvzV1F5
1VFdGG1x1mf7B6wLkSf22A3hsVkBCDF50xtUegwvyMSrUUj/BMulH4G0zhUKTynJQZSCAW7jkEOU
6PU7SEF6wmeHaDliHav2UTcok7AxsqTF4vPhU5Cg40aEQYBRxFMqVugXlzRW/aqcdHQ+128pmwej
dnVuZ3NwZd4jCiz9Owf9t6XfU3LjjJ5Gpev1DAUjn1d8W1dn0RojAEQsGVjwPcW23UTSayn6djEt
EvR7vp/mqH0OwH/k+U1DqreCtjAMH6XSptmOhSHw88Y0+t59VFz/TWJba9XseVg+5NEsgfymvuqW
+phZJUUKHTnIYajhvFZn7POmhmRT08zKIzdeZ4EHIg6UbBhczAKIS3B4ERXUvcaGlshsL801fhN5
7D+rFHq/cNpVi3j/XjCj05XZjH2Agp54CTbK4wY5DG/nsmMDtOspd+avtC7Mc8uq60dW31YEJT5l
CtP0gLObqGPm2OGGzSpLtmdmIRjLEh+DNECgI7bHWAwhxFZYJ4EQjvFFU9xv5VC6NzGGIvQzGvxl
J5bd81DVlipdmgaQ60pODLGKbM3B4kRTHcdWvvFrZgyJ3d4uaYLr4Fs6qSk6jQQAU7p+IP9hViun
AAxAFLVAvzslgoYWSDSzniZ+UrMPmfMwwznuX3xA/xFZ9ZsEMSjm922OwMhJ6uDUUAEgeFTNk+NJ
fxm515MPM6fxbBen34CXevczFovpyfCjfIkpy3qfzrlyOJOsNskxBsde/um/fZdcSSsMpFltTDRX
1rHZHyt4U5w5npfSh2EFNI2ptbe8/+kREPoVcYDSncPU7YfmCq8SjgNw5mlVnbsyknNckaQ1b06l
mqZBO4IIP/EHewCU5rIa4KY2RXPDxYt9tZMxKD/zOX6T/6aRrKP12fuCOiGuCEZsYFfB1qmL0pmF
U/ukxnxFEgM49SUNE9GyMZ42FiagQPNCwsi40xsdnxV1ZSr4bw33D/M4c90sRUqFDESViVxHqgO7
Z9LsVtF16I5KpfiowlGELKjZHyXN/oQjcIsbB11AZEnOVxAiM0wTONcdfHDm10HInjTcATQvbuOM
j9mrZcMzAKPuIknIRsvDqff9fttnQUTOWx+9lri5S28iuscE36/Mwgz32fbw1IkOWnTtvQD9BdpE
HHGx3eg+RKEvCI78zeXM/2xoMDNmHJgsJpJdRa5G3vgXMETqJI85Xtc0usgiWEQaWJkOHEr7ZDTJ
241marL+68un5l/dWaj24kWVzFFHdRlVKlVnC/+3pVCmTxbfh5Sa04JagT3K9+/kuF06Un6yAMjb
UnA+cutxUx77VN8ayFTpPDwUiRhEhXkzvuSuBXKLIfUA35Y9/gghpkcloGaD+teBgaNvKarYacYZ
7IFtS+SqbDFD4tygL6E30IRIGKg8NMWlJaZ7ujXLjQ7Uahm+D+mD6fLTAHFcORrsb28SN6//mK4g
NyGbNk+HvEltRcLnmocg+KEz/xGNqr1LxEV6dWOdlKMx1EkShHqM7gK2QhF38M35hWmq9DRl21MG
9RWTX9nEUpU6CkBnmyabQhHS268iYc3nRJ4OrEvnqI5RWsgI+T64WSkOGqa23YnN3HneaKMZU4pk
qy8FeoxOXUP7z8NU+jeiX7FNGi0lPcbn7A1TfkwSFKbwtM165Trvb56nw6Jnd/I63jmOEtvwQiSB
AdRzPVLt8nOx4CSBZWvA5wKGo5C9MvlsxmpXC93lyXd1PQ56t1t/y0PxtGqoSazsxBExHp80Mo4p
S7zXKyYenOLIbH8ZpE7wSSIYzltr1+DUwz3oF6rIofdYOgDGF45DLfDTRbyLHAqZET3mzJuIuvkp
Eadw19vq52ajvXc5z4d6jtrkOfGkv8O5Se/HQyD0TAZNObWnQ4W7XFOafNVFlkJNG6xt9tgFAAQq
ong4jYTzKl0Ei/9oa14GK+IXMU/N/I3H9eMblcxV6Vcgye94aSOr4rZx43RniGTjabGx5Ef497m6
Xps1VXMhp+f638gUR+fXFSvIQp1h//YJGiVnHVATMGK89G0axthfDVF0+2L2oQSu8nu2yxD4du/L
1RESEIMH8aKSfWr/vrU9bSdKn1cyoXN1Qc9hmcYLaXspEZdzuTFGcaGJdG4mTOD5wYYgA6ooAO4E
CPEosKQXTxWW0D/P65LvjRbH5rsBIeNlnKv350YKVmyb9a61n1veq7b/Ha14CxbGaFXRalETia1V
1TiPSilze6Zof9v6eCIDmP3vCpXM+k1I4J31ODfAVZIcndewRONJm+ZaC+H6ISz6igcwjm8ANSNe
8vbuQP37oJdBN9+zcBP8mhiELLpuKj544ivZbJNruoE5FlK8qkB2o3EwqMvBCxwTTZITTEWctMfU
r4ZWkkCrRfT4rmUvU4AutczZN2FCNqp4K5XEmEUlN0mlYTq1zHy6yyw5Nb5PrUkqXACsDL8mGDpE
As8IJ6+DNw45xHs8PEXGE4YMJ7OJO6eKQPh10Czkt7brJuc0NxTv85uf1yGi9m/6Xeuhz99HiLe/
lRH2aSfPffzMur4LoakYdkPk7XmR3oKpAT46O1tiFKs1xR23x/+14AXz+kQlkN3QZKRDBx/VKd+v
p+TllXX/QvUiLpgK3N8Q32RnC5m9mrCOouK8JYO3O+tFbWatvyChm5eqkECaex+Cajn6JhshMrXe
lOuyMAnzT9g0y9HJkurXgD7TFSO4KiWHQkzuqo99e7anCn+zM7+0kXMbNai2f5jq84fgjYRYZ6xm
PXTenA0SrNyCBsevVIpURLK3HN/lwIDlqhuJZc7vcNlwqE47m3EX81BPsa5H7tep1hOGDqcivvmR
yhDo7+MJOIacnLkXVW4tOacgmEj+7Rn1ZxWmPFlyJ8qQlh0OaEiXosYW5m4zY5LITmQdZNkpjyAz
T1IVXbmts9PlXlR+5DSsLAUJDoqep4VbPaI9C+Zc0MLizLspQLyI/i/ZgX+Q0apIDcNhoHc8F6+h
vdgsP22QawkPmYaLZiMsT3kpjYW4Tv2q1TDR19UfhFsl8y7N28TkB03Cf2L/uA5lYbOLuJYWO7D9
KkhP+dK/BCT0pna0UOMxsldcoR10hjC8am61g2PTjZQFnYmS8eUBWMgz+fIvAx/h0qq0u5yIt/1n
EsfsqU3hurgWfvNUzfU447t9yx1PJCdMGy2Y9e1QmqOtTZwVwBK3u1I8T6eUXx1oQ4SpYXTOCou9
F4YawRyim1gDchc5RTLSwjVhz0cZJu3tsskxaCMYxCPjs0aAMHkABa7pzxg6OdgtvQWVVEUt70Md
N9Ed/VDxJsimln5cyuBEO0aggImgiSbgthHNbpNLCYMmBjbV2XiaULP4g84kGRyJlSh5LD4E1uLP
eAitZCUTUs/4s752Wq2P0oQXK3o74NaRqsgpnkdLx43uUR8V41ZPDnwFMgLhCg57b9aHQVYu8zu+
tHTbAOCFfIqU+W2CPzEby/sOplAeDtlvaSGDr8O/GyFIgwd78SDjHWLhBPJ777Ovuc6ezVb/CKPL
5QhFFkS0VRgy4PAE0MrD2VmO9annP5ZDLj+fzdc/jmwOfZff9UqMap1C/tgPrYLNGXjX/qW7kTLv
XDmYyZwusmc1DrsVZVpZU4zzK+jw5EuVieaNgC+Ic02fGD834nPoDliB7nkO+9LF+XM1eiOS4AFI
hNm3Xpq+EVfDbeBxHdK9VdDsZtpOcxNLZS2ZpKGK9mbEM2xgm+wPP5fXRmeyw+MUlDiU/nh3/gz+
K4Bm/GQiI2Lx/IKM+WUUY+dMl1UgT6S6eOLm6NKXniw9j7TXDWxlubiPakAfbW5XMD1ZcEha2tdK
TOdna/5YW4BAK3RoZTfgPww+Po/sAMR7nEuX61cwgEF2tiEiDJSgbUofymztTQ00893tvZtF7+rI
SeoPKarPIMHgqPPwDYVaUjlxI8bJBtcClTU3fkN80OVrMc0HD0KxkyJrZVYHzdQ2e6HIhdYaSYyo
wTshyIdL0mXGKD/ZwckCQnM7PKv1Kfk3tTQdp7qG3D5PnFG9daYadlR1rN0BKz6XCgrMPTCF72PA
ZNC8+j4tXtRMP4TRo8bBI0xT7MCN705OQURAjfOvfBjr7kLyQWmHnWEXFUSl5fSfKhh2RMvFKzQK
44CZQ+y8L2ZJpJCvLmsgriLGMZtqMAokOdL44D6B+ZPzR6reSGpxhSbv/hAJPjdd1VzuK0JmkYLD
uZ5D/a9nWX+PRSu/E68r4xmP/6rkmlWx4lC01h6Ol+tR9v1NP3VEDj2OssM7uuPspAHyB1JVvojt
kMD9HPySlN9sGK08PxCi0ByV4z7gT6b1jf2WScN5BMI18Q67YkjkuhLigusTZmUGvoKoTrd1/FEr
gOUWCJ6zsEmPEtJQyhCdQgfZTiQYLYqUMxn27DO6BLDT+SgEVI9rmx+lJFOR0WJWEV45+mkqUDtH
uJiE8p68PsARfcqNzZkvnESn9+Mk62vfz5zkHSlatJe4bRvMcN/5nG/PrvZK4mXUgrdH3qh4nTrl
mWh+2N/ruPWThls7OgUTan73Ce/cThn+ds0gL55dOAyCqCBHrMJhzP9H1uor5PXiJpZMoVSHH4w2
SRgsNiftsXC0mWKCTkhc+hqRf7mzcyTZi3H9JXc1pWurnwmYySkzBLewuClXq3AHZQOD1VCsz4Le
D/QbXmWNjs1cWymjKilLJj0YjT3eN/SzS3il0ujpuLEZu4eGdaS0L+XXGACZJ9X+Boy43zKUQBUG
dwIud2GAYJFwvI8a44oe3lIRf2nvC96oEu1plnaeTgDBLuEHmG9EoWYg1VZas+okeFLWCwJyOiar
6afff/R0KCWr8f4Gug34x1VUkmxttRLpMfgybVnRlOKzDDTaTgIR0++VrqPv+dxKTB+hmU5dqus1
YPpnvlfKk/jkKQ2lU/Ln5TVp+jkQBMPC9SI6uS75ZLGCQB5Fac9pBDBHtg7E960fk6goLgCIUoF0
wpn3Jjg7Mkj3VNjeyYtfBDp7+F2bu3Hvm4QoDesVnM0ULhlEOth8JgHffCM3Ik6k5LGygIhnCo9L
HbGnSV7k46/rctw7j/eUV/j/ZnK8FJY+3uIf8i9oFMQXz7ERxrRR9fd9NTMZnjFRi07sWgNhv5yy
oHUgGNTRk8h8UM5kFxhKLW02RlcD0W3PnJ7wtZiiSnqCvSVXDWWLMBxYeuvniuWreS5Wp0t5pPuN
fJo4rD1XKGTEjPmFYgYiNuy9r2jKi9nDesu/R8s3O1Sp2QiA1Q3d8X91nj4ZchXMTbECEe1kL4OO
gICRlN0rEIqMG8l7O5WQ4BCyVd1aQR9PWKpiU0tWMAErpZ0V1OleukLxh47PBYPtHvyhQqIOaFyx
dEC1VpQV6HTHFbQF+vcHvNsMu4hoTfHzrvaBZ+Z847wfhGwFPrTxaZMBggH5QpeQdZ26cBIJP0NO
swW/loNlu2cRIJotQOJu+G1Awu5oY67GA+A74cIddmZUm55xUOWnhKKJocwAKf2n9ERQoZH26FU9
QTpBBQ06EBY5HAXfbns+SjKJCOcv7BMOJzez7N9idco3Lof2GtPgdCLyWTxJXI96xEP27n4e5ujI
Clw2XUxn7fQ2vUEk/wNbDJ/z1QdQfVv7h6ssUkxVls5Xdo9iQ6ywbqzjAyUOSbRYYw+kybD+4jJI
qObTVnWzx2MBSAiFXpnzppCncbgzS3apMvTqP/PQxAarKKhE3amWljZv5FCLSnQHYYdsI/1MM2ys
44V1XkZ6suwScSzvLh6HFOI1L5YpvZVVINPv7kK/wiodraVoWh5Rfgcz52oQ96nlpSZyJ2E4BIlZ
kJE816I4C57HuVzZPkWPKlbMufz+1vBYtEq0PGhmQQMvbt73LaN147TP/6s1KrRfg/qgDFBa0OED
KCGlqRD2pq63MmQ6n9LcR6uSc37nyn/zZ8NEMttK7tv8W7l9bqwPWzD5Vh2cPaAsJwKZfhmLxVU6
p+Sy86AGgXfwQC6v7z2qLQg2iPT8aeNtJqnvNqyBfQINRuOzoDzvyG4BRAyAfNEPpXaFsMVDyVHa
HdkLcnRSAjg0DvXzOV4ELAjiP8kMg2nhzgSugQy+6hOxvwS/6kdVJQO7tCWO8FlNo0C4M5czjm5W
icM9GcuZfOcl33LgKkysMfuF3eEyNYtATnH95nmK1NEFBHnfSKoDDeXQvmeGzU1qrzDWiRCfvST2
EhHZTlQP1R2CCFLuaaSm9F8+NPG/5XvBTdu6sCeH3MEzAQmNFV8seA4vO4seflEYdWTvJw9jDmJ6
zIDJj5wgBkzoCaOfosmYNzAd7lnQJitz/+DlFWZ4U6sn3ywP0FbFfTRsf02fcM5ZbczeCpcDAl2C
sD4ViWMRPFcyfGGZZmTMzXqGNlq5ie8Q0x+dJV1JfwbvdrF8/Z4PxtT58fAbUt+cfLBYkEv5Bb0c
Jzy1pZXzSLOtcCB0LcTzLgz6wKCDoRR0SWC5nDSjU5bNYxV4hGRe5hdQ+KbH7smiSIhFkeRPdLjR
cFRsH4Zr2/wS3kxs7NYeanW8wy8p9twRSvdqxVBCq+F6K/JgRobQZl6DWdIA/huR3YpRS3n09V5O
GJoxhQFsNBbjo1maGvclGHf0dTvRDxuW4JSHzdl0zR4ZWMRTVzINaRCewVQdZgLVZ4iOV5W0h7pk
kv99F41EHwd+BZEtt4DpZN+903jXJtC5S2Ox2m8D7BaIO5Q+zdqyhWptG7x1kzY261TuEwRvu+qB
L7FNSEIA6Dd9ycIL7QOqS1uecTSdsj41iigWqOvF1EaMWv4aiXFU8T+FqIrS+OhPE8LtDrur6GFA
lXKkHJojNarfSK1501DJQ1N1GDPExYEs936sc/OR0zMIPP5b7qP5qHVe8ot7mzlRfdsAjgcg5YhL
Z1I+7s28DfL8lxkkohYuTVgAhTX+ItIr/xR3m5oaroKYdJBk5jRfrcx1rfqdLpxxwvz964gKGJ9T
2iBRitTo899Xr6Tt9XwfOPmVEoMfGLrGc/awEiJVN0ZWEnrpK2fhjnWOL0plemsivD26RLzGR++q
3qCUU0JARjSn7UGo+6GutkI1ol0+MumHd4/QpjXtnOtJySAzfX8wZP9iiQpGoL9RbxFWhN16db5k
ThITUcO9zNPvFObx+qC8NI8e3ChofRu62ZA2ZC9mkJskxPPFsQWeSMA4Xa0y+ieWEqGjAd/zbYLA
cs/+4MYeQpObJZYDtRouGp+ilWoheePLuq61NY86klHWy69XnFtTPDyUbCwnQGnjnGAK7wyy2Gzg
a69lBbAVgnNAPJLq6PP2i3p0nHmPNQElX0lZXm7eYD1F3qK+1nA95/DRf723oJOFj7fNKrCliWj1
KjVWfwoa9JaLPcTx5IC9/09+GhpCa6BR8dPk56jt5l1nTCUaXtt+IwdlMx/kddh8rLNhjdXoVBam
OO8OIAsEiCypB0k+pIyvIFKxO/vuMJqK/n9axYjj6fJEXXQJXKrsbX2uiOrUgziFK6SGVcVIv1yq
NjBfbrGyQQ29pRAxzNBWmDAQaXqtTSCqOncqJdOfiKbTri+xa+ZEop4KbsnpWFt0d4gBCqnAxix0
c7+pVhkGaqAxuFiXTZPYbwxLYjUE+NL5mrQ2iKJzwSjvm+vKdRADppal4rHa8GIE3OIQYdXosAdz
sekaxovv36dWFx5LEj1uRpu0CKcC2AwDf/pHotL8oQLSjIBljWFUY8PNxZVQsrdPOAaaL+JjX6xC
mHYGm2qWU/rVU27NNayOkfdaVpQgQT5OLUvQy/VhX7jOIw/kATcbdhROZfVdMALoyN2tnT7bptPP
29ra09QNaMU+9pGkD3+5VT1hR8vWpoExUM/16LTxMTfj0lFZZgaDRfgRRb7XBolvG/xUAgvFJpy8
ygTUJjUQ+A6tbBOpCFPAHCpxLez+zvBjQ3B4bzaXZ2KxnOVsb4jVeg1hoLyd9YYxYRmXwujDUAip
8zr5D/oSA6HWIx5N52ZTLOiq59SSFSPHNYsMXjc95h16qiQy6vimjhZU7fDDZE9xSjjK4odligZD
yHqOQT6KYEW3kbuJz4Pg5Jo38cfgyzFuA6Y+TRorR4X6BzVLUrEKbh6zSxpmrfYdIgTN6lz9+8Gg
Ro3/h3/uPM1ZyucCt/Y8nXgtWXJixSdKuTUUgSyfScNHKHhmD6eap/DWKWyAKbw56Raq/NfXw1Lc
c0qSJzUsL1sLk7ZxFPzh/Dmi8WMcTaGlNgCZ8ESwrAUeeYwHfHmAY5xWaH/B+26uwb0iGhoNv65v
FE3sUdE2ZtgsElDW0AM7MX4Uwnh9FsIkljFAIgPPPpLy/znOKItMDx98hu2ndv75tKYkK4zJEQ+m
w+pBO1AYq5xxNvNi7fLdXwM2QCF9y4U2anEtKDvs5jTJ7/2ZjCk8sf4+qCGkIY5JBpXyLNpRyL6s
+m/bXQ4xbG1V5JLU20/esZmwjrct+y9+W2jShHy9UNaekpRUW8dwPbyQ64PhkW60YHyPbT76yV2W
FY0RxEruuDMh+6dWBoPeuATjUBnBhcJMEsEe6qAymwCZ2sVOXwBa2jZrHAC5EIhC+9c9SkqwCrWH
gWYJpOWnE9lYVDjpszpaah7SjDEZrikD7AnHQN2SKCH7U/ULis+rVgZTW9BmwyGUnCpF7Xxp8iud
XmXnA68WKviJNuq670bIPOa6Kain3econsCH3Sm0KCp0hftJawOMyNigHC51w9Rk9GB8p1aejxeM
6W2LAzxc0AX1d6lW9JSWlXkCClNGeXkGwg9Q0DkSiKOp4hJ5ma4TWT5E4SV4XslHauk3BXfsILzp
c1/8FyC8s/CXNTp3/TKh8TqmCecTOCO/XH3Atwto0QocXVvCdFprESDluCPlo4eweuU6/PtYsf8M
kUnC1PJqU45SUxoq6nBsmFOlYN5/lKX3JmleCZK8hKKY7NZXGFVNevGFAj7dvIG318OZed9rPgMi
+pKWaEvmhZzi3vXY4Wxi8jibqitrifunG99Bixs3ckFqAD23yDnDFrZ/jjXq1KADzKKr4src6YBD
vzgzhWM7WSE202AaEMnZF6myL/wxBV20a2pTBe+dYx1xZFIX3Nq9PIuy56x8ejIIbVD5sY1NQ4uA
neaSmXgJs8NQ0vfgz1ZnjbVN6n6mGsGmK4hXpB+U50Gu86PfOmraKSVHLZCd3EtecEvcs+gses7m
kNUk/Iu5WafiYr0EjW0hgJTHUCvDE//rmLVAO/a1dVyJbcoePGwkL03L2J2kD5EZaE+S6CYbp8fw
JXEw9QMNxYybgPdyxP7HC4tWpATSb/w+uZKvvShcuXelXv9c49R/Y+8HZPMxcJ7zK+wo2o4EdSW1
Ucg2GN1R5fdBQSeCHkxn6N5VE5oyjrBgqp/RxdhAA105M8NaAcEVLinDQJ8CCFZkm2aThpejVfBH
CeaR8vtXtkMeGXwrel1QDGCJgnCrmY/EvJbCtS7Sbjf0OCX8YyKBCu26nhp/gGTMc0RtHzQr6KVy
iAXZcWzZ9XTAnlcAtHPcnFU4ZADXnnQ+vtywiA+pYkWt1cID0wSqV8A9/nQWkxbpzBtK0q1Qc0p9
pliLO2w333vZd/iwzfdGTKLoen/BUnGJWwEzNkI79nSyDVHwQgwYrtFHL2NrYcbXgR+RqXG7EM1c
Rpbi28lQPHUlqB6+t7nX290LbHROCIJ4G8Wts+W6TBa6NkpXLHWYQ+L+WGNMUwjddmScNz1X4PGM
CMDngJA9fx9UHSAUxcbT9lxGtwSu3ri5308fyhR4B2Q4htt3Qr2f2Gmycx5m/kf6GSH0fARD4QNd
43nf+TMp8QSkpUwMd79J61KPZAkqoLRLTxrLs1tJ3NVsJRzDQfAD/oJ+sj8SSXn/SkRnBiDO7vNW
Xbnny4j2tO/nSAK6k7bB+TitGImXzuvMEgfHXcBj18lxJO6qqVjzQj9cQX0SebZfsKWexmLML4nn
wugUaPrHX0Tv4ZQPRWx7vemNFxMoFLEUe1io4VvFCXuw/AM+dgJ6rQRLStg3CCs2hAdnDBXu4cSA
gp4Q3fwI1Vw4P6RqvTea+DWeuG5NH6FFEfdez3Zg81wU6kOZw85/221DahwafTYHbMEdeyKzB2Nx
bnr5YeVNcxsUAEMB9e/hlqGPFrBcjbzmmrnH6D422o4qIwMPPQzzCtJOZDNQjsl4Lb9ACjg+tnLh
LnheovtiNHIdZ6UnZXig3wilRTadhAedY1EN7CNo+dV09ym0P9zEPUSjTLFkA1czse3jX2ajVBaq
2loUdchlXK2coneK44zl1d8x/svV3lqMszju35BvEiwuM4qdSnV5DGaSyCPyJJ7O8qL5jmfYON3h
erbxqhtVJp0uEZ3YprQ3XoysNEyC/VOoCh4W117ejhwe4dGSwxJ2cbJtu9n6HPf0CX1GYriLNZ4v
8H8z58OmTRQz55UaKug8ckHmZTnBw1fEg5OIcQ2xt9lFPNCUJr8FJmXQ6MjFq3oND95lQ+p2aKfE
3rVzEVD7pOsCVs3rNKsKvpEU5/O+KNABO3/3lCvGBeJPkXfs2qN3DGZc359IAnnYM8yJ08Ha2lY3
EG4uwqe3G9FztrFv/Kv0jHsWlv88QLvX6t5Otc2BToKpOIk0oPc9pBhj2MmAqFDCSIJqsGIVSf3h
hhIrozlNHJdP7srQO8Kv9PCq83ZWk9Lz+ZcuQcvHX1Q1mNrz1bhKpLP9jE+rkkczL4tV+oldsUrT
UR1KcpvWNFQ5al6qihJwYDPh9bXq/W2eXjyi/lSvU3LK2HvgGq4G3F2KRndsyZv4PgDIBitH/LBU
y1gyxqJNTZg3/zGnIWnFe1w8OEAM6yc9X5ZrOQr2WjicvX5eEVgetKWkAzjCW3c3gamDQBnBC8i2
Z/5PGF/yDfhbHy/6NSh/60QBFht/kUwhXuC1MhbGGxczlq0IZ4qIk1DtvoGh34Ri9CoXRXSb8h+Y
Ro+rG2PDAwlWhp0u4vNu0HIZSVxf02DaLYWyX6ibbhmE0KsrOfLxY4LX2sLKleC5vYHoc2oYX6pa
hSiIpc45piR8uR+qkT3RA+DbA+jdTUzL0NFUtUcPapfDb9fwvH669cqkIiA/GRGRoBWgklxlFMHK
i51u3H+gaku5U2I3JMQkVIFXXrLq4p0xKg0VFU1i4pZUm5HhsWluXD2JKe09uioKB09+b3CySNBZ
YEBlKnSduTJu59vsuF168Nv3CZRML11PizBkOnSri5Dkz0vVcBuHULMH0r1ToKLJvOZyW47KGZOR
vYE6l0VXMHlOHFGTvyFXoRMlaH8HoxJbo4uJNJQBFu9khXrmWCtQUjTujoVLcbav7m8yhXN5ezah
6tSs9rrsxPyfMtSoAipKJCBVb0dutlP+fXqypGi/nometEuZQMeNEMTPi27039p22AIcatBcBsf7
OFGONad53pywoUiDxtybf0h2l/6PxNmcXi87oAwlGVMfiHFxAWnz4tLPms+Shs2ftu2p+/5jNx5K
psjxgSTBvPjz/Qh1WB3zv3KN12gHfUwLjdsL56uOvKJHzxhZwDlgmlS2i9vA7xpk0I2UcjiV75ki
BDW6iXpcwxtfZ95YsgVi4kkJLh4fntZuhBuuTUtT0bBMXHujlJVZTiJDP1cT1QNeHWilJSsyHpcc
SJGcWvhf7529Cvzvlp1A6BWneVMzolZH62W7V1gDF40t0WGivuBbh70Vuxf64yvfaxbqLGNB6EPa
YPrX0CqeXm2YAt8ZEdn5M/kzBdO0Qc4/FjBUhYB7egLWziRk54v+CdyyNPZWpi9TDjY/UtCgqlwL
x1Pt6PNZyWj7h3EIMt7H6/FInAZuW0b4VpaPAVhxmvjmOvSPwV/YChMrTCQryrauNcSALiGOnwIP
dedqKqOw/x2dJUyzjS2jcYTWN1OBnU6SW4JUV8soHOVRj17IbAFsW2akH2z9CJ2RfYsd9fx9sHQC
TH5QZkeqDY2DoYZyljTfIcBv9dj0mSoVcYfnnfTRuGfu51CNKikMFSmXSqU3vu2BjokEH2kp4KEk
qrJGhq2Fj1mfsKoc33JWQ0nTy8VmWxUhyZUGCtPul3MZQSi0/+PJMnnFnbcc65TFC6flkhRQYXFm
PQGToj7Sw+To1ecwm1j8WHHLHo33+mRMPgMuEB0h6ze3fHxkjeWHIIyODshix/vyA9BvibQL//ME
xercl6A9mdx1ybpS//oCUYFedCTvTGz7gw1FGnKfOrkSsbpqobzx/xGIsLnR2E/wN/ffTVp8T1HN
2J6HCXCv8xneYxK7bR+vbDEhA7bYjK7y5JJD7ZhtiSJOfRgr6J4IIktA9jXYbxGx49oXzZgUuQLt
rEqp0Fh1RRYGw5209xYt/36Jt4gcJFIL2PE3f+Lwd9YJ3wMtkGK1BVCgW1Hl49BvU8xx5OBzaMBE
sS3TvubzKsyicL1xyJXs9jNAIwqLKLlzo7u1765E+QcekPn2hcSqSxhEw9xD1mxklToa5YCMOghw
JH5xuAiMBbxAGaODqtLV7mOWyoBP7geTmte1UdYpJM2HWoFrZs/wamP/FL4Ax4hi3SAeYCEKZ92s
s9Mx9AUnvz1HCAhVdehEWnxX/Xy3bQr4Ue4Wingicrl132Aq8nAS1mPU7LChTZQ2rHdFcqwJkflY
7k2x6jKyjD0uzLDH5UdRI+yENgR6ebH/nMImeaaDlPrnhzXULMHS+82GqVSuW1sFnIOBa5QIs8cx
BUYZ4dmFH2SMgUlr25SHPsAJC3NNFMOx5v2l1vbxnWMFGZ+tVu5Q3cfXMkCADnIvA2toGm1xT+MY
VH4nwLX4ESn8kcn11ZOf3oAU/suWK+0PscpPARsGGnVyYtumAMwr27Na9WuUtW98bNglpJ9lkm2f
9Qzw1FCsV7UaepgngNG0ZfG3SjqP8M8uDBjvvGf3uHJYGEV1mk/8tPBYhtz1OpkE22/iK76Mv/wp
+hXpWflLj/xHvCiy47pYvrhCzoIJcNbFNbrYWHkNqqFevTXi8lbVFR44oCC0P9A+oCD5Dg6ykq1R
d0DdvHwcKDlI73KSXVQRPy+UCB+Z7cslx83LsuRkss7QwZBhc4KmQwZ0aYLyFNFhzAFvY9rhTUFF
DZYxiMAK3VY6HPoPBFPSl+PE1y8OW0kU96ZRKi5JHI/DuzdGf80mhzTcnf2ayz19g1ls18RFrTpl
5/yRUt+NQEXhpcQMNQ19rwOnkj0cnGLq9q1JDG25Fu1t2iwrBAHe3ONXC+3lVZy6DOUhSD0wLc4O
YYdfE3uvLjPjh18OY1kckQ62tHC00t0wH5jJPE8lkYOLnu1K/lYQcxgQLg1m5jRJCro2ec9Loe3h
hVpn+TSZDGs/K06umMfOFAN3SIJlX/QRjowyuMTpBlcUIn+BuRUlxdXxPl4yMNOrV02Joqzr4Sm/
IVVKPx5aBCekJXzKVdHn4ZJ5+txK+X0jsA5iiJ6ILnCueYPOHLkfB+1MG/yKOxk0oVeuMDdHAedV
RPshdZtz+O8uGRTmihrCYr874FtJ4PAj2J6YmOE2+wrb9+35Sr++P9fOrcrZLe+mNi3tPVyWw1eZ
FlB5U8vjzYyttDJqK1JvxzxTVu9nugV9N7DAEFIAbQpBlSNvHynHsTSa3Pf1GWXiYZp+QLgg/Mer
Gf5dEcaeSCf/LlZzzq6Yu1C2y49Nr/D2wjJsrFSneIZDReYhnZoswMQ5KxRBwql4B/ubAGbh5n1k
96Qi4kI4TZkkf/MNoGY7MIc5ZAboKlWGcOKdoGY+QwiOP65XP06lpwwSpGUj7EivTMrXBfQ2a4r2
epscV5m4gnBHqU59MpwQrVLK3goJx9da5r0AipRUcyjYfN/Bqfu/MtW/3k+JF7v44HQq3ht+BuX/
w32jjWEh5TmPiICido41B1UhtmzL/PcFKQpIowQgVJcbLnnqI7z6dhzUaChXH1EQQy3xxEQj28KR
QMvCbPEEFunPbOPNCPnybu1gm/dy/0g6p+aPJ8uFldEoiWqCxKEIb4DjC5cJmihuf8IvquKc34WX
0JP9yeY8rlvvFxcchHJCEb0GARkj51zMVlyF0s0Hc1q7fAeiZIQOJ8r+GiFEptBMmIxnn4a0K+Aa
KLDmjfNItmM9xPwY6UD8MxmGuDmmXM50RlGg7M8pPYiuWWMzhlwTdvKpNmHI8gD6d6PIZ8X2OXtE
U71ZEjVLoLA7IHEM+wG/wlqo9ZHmGa8WFRSDS71qyD4QTCKlLgfPeMnJjFp5yVoFm84qW8XuZWkv
SkmlxBqla2wTZUc747EH/jP1FxDxzXJ8t7EVe3CaQTdUdPBA4va+6JiZ8l1tRFZWtjgHIbgaWodL
HvRFHsjGf5oITs5xd1etbcfJr7HX5ejWBXXAnL1nxEMh9yVGllJuRtZHErfx6l6QbjxXdQj7k+BU
sQCnsj6/BIxxeNarvHo3pjR5BF+BOgsiaTM04dLEMiQGdV+mHQlQnPU3a3aEnhoBmJpLI6gotusZ
JPoaSyYFf7j1/XObJFqH+8ha8i4tzULMilaXktgEQ7jg1aLd2C85oMA+H9oYAWAgID+pKZ3SRlOJ
Wp/nT3E5Zc7+D0xpXlfoS1y9fz+ejusaDcbrjbq13oJaZ8sze7ynGM79lRvDH2hnlJNcQYeEU0VV
vDW59MYxGTUBzNC5b6BDtMXwTnqKA7dkiaQ2qjRbsakfpC20O9N8RyUGjFGCyyhOwxnXB8BrQER4
xabb9PLI5+UiKYv+d6HYkqNxUweb8LhqL7/PrZiQ+qY8j4U7BTvVaV+5jsJoXxVMtjKnvj9kxByf
8g3W2qK66TPOeajl5sIec0vTxrt33V8eQkfukPw/5cYg2RPsRHvHQqKL7tN2RKPu4JGLJ4tVSwBE
lUUB1p0DAC4hty3egvb6AUol0T0c0jqfpnBhjOIxK+6g6WD13gCrn9l661tVSB1IVTtByzcoFJEy
/SxlT1xhpSIYxf5O1vQfjJbOasTPykaNnPMK96JrNSyvO8hs7hx78fRIVdQemIDNE8poB7DHChcN
zt2wvAPT70YKO2tA//Dy84WlHK7/TksWz/psSmjz0WADHRUZK1JN6ISWX0khFaLrB3Ip6NJja1U9
2L7X/vwPRQKV65HcVmZNCrFfV1TUfm9zDUq5O2Z7Xakp+j0dRpc/KGOAFG6oHf4Rx7TmQ9kperU6
V0SW+W1qAlY98LNsLcLtdUZK7LOxXu+Hp9mTMEEEXPWfI1ew/J+KsfmOjURYHunbGH9nPG61jLd8
yH3/9Gz1+JYRU4I8h8nvAh7OQYbHBgZlv8ckQG6uPXmp8znvDX1PLT95kD2wS4hEIqgT7xbxa8aI
IW7OwAS0GrnFdonQ17AayIsMC8Y8RYN6gg1asILF7syEsi3IeeITexh5xDhMUOlwlLi8fMiwuLfS
XR5Zt258bkAzAcx3KLjyKQ/zS6J2KubeA+uQe3GBFMFYoVrb11DeVmhRTahWjH2R1Bui0162KxsT
CqZSgCE5jf1uHUH28FDcQm/LF3oRb28NqJrJXAgIJZTLqAluJr3SBM1ScPbDo0T2SG7uxiYZXVll
Kcfsqp7o7+DzJRQr23ss8QjEfnzk1jKoJ6aFBaYr339QUdm9vT18d5Oynxx48euZ4a0YO8xBvL5j
0KcQwVTL1gEE7bBvUwInJCnF8/EhnjxueMKlYLN1hhDG2h02fBpLDUNI5omLhilFW4BN8FQ5aHdO
PNLrNnF4g5dm864f+Hz4/AOngMqcCcfZhTQ/y0kGgiH4J/ufnHRub4qFwCfVqPg5kL4/WxztW3T/
rHmh2/hZLrlHqC6BGmsY4SCQqcsJfkEkzznfuQmGx+JGKdI3ac+3vsWncBNF9M6jN0uMNxDTxOLj
4suZdRvFyvFQtPAmtEj0QLcuD6UAg9IMu2scwm0eAw2dtgNg2hiS3xaYyls8c3CpuzY2wc2drcKe
b5Cl3CjR9cmPDvm4DRcrtYcu8lwDOS1Dl7E5jFPhrzgUjTC9/9gKS/WGLeGXu45dI92OIM9NRAjI
r1JSPWZkSptRsD16DYiwiB6rQgj5Onuo01AHD8+fE0e8BeRUPpyyPHU+YfSa7uEeQIUyBWWHw3Qc
eHHNyLSypTQjVhFvwSJjpvq48PvDLWpCUISYI6AnRZy4gla1tEJtVuDi6aj3vX+6H7g7qxzTKwmS
TKiGSO6B9ihdJIBnx/yKm8wyc3KUkDbkQaNgv1coQ6wcNtNrTs9n94XcZiowwQ+j2husYYkK7Roz
irFUApI7kw+ly9geMl92jsXPUpmvJrpdp+RemLBhlQC5Ba28eRZhLOy54bvJB3VzdieDLwlVeD+g
XDxxz5nl45PpS17t/mHBGiVQZIv9x7LlLN66SjWJJXXOWx214mmvESQhZh8mM+dirUJoMD408Txe
QHsKQUfoVVh/YbpppCbQGAffZbnwhzDMxXOkZiJiaolBTVoqE2HeoO7IxEOlVFDsNvyMpykCSfvi
JMG20ul3nFZl3QdH8q2v9++eaEfZ+q/PW6zXkdWGwIHNgpRl+CyCmMh737gMN+Xm7R9zQdMAo3tn
JZYLXXYe5YmJ5Qiur2zkvk3DCkbHDbqObLvS94h0PUdUSEDS4klYvIC+NhMAPFCHm8Z6kWYiH1ua
IBWzmhi2WGd3ajkalfCWRVYC1lVF7Sdq7u4WhHWSntCHOWxIvvgtsxec0x2b0Eu+UqSk2ydAMzwI
3SUWZvc/+SKTFIcV8RcGy+OzCjmVQtIwHj5GBSrQw/z0FcEdvbeOv5LLl02pApdo0IUUUgIJwZgX
DmzbXas7pGo+qJGlyQgVgrP5z3em5fcdXydz0y6KFg2sVQZsh3qIivwOr6YdxtL0pYhX30+xwiPs
Xqp/TWq96xQV/253IKuMT2SZ5gnUXM0hUMQt3IALRe2lriGyF6JcMCqBJiapkcZO0UxVqtGW20hB
M9FfFt8kkl0obSp5oVoz14wQ5Obq6+Bz89nrYJCkzH1ZbhkKEgezoez9wlhvwIoYmMSER0Cp48jN
dGgxoRuQMHczhPvVke2qRKpS/TgQ2R/Njmeq9DJ4B/SKOxhbf5bzrczMGJgFxA+3H5XQjadIDK/r
TQoQ0+KKb9g43Vo9eowNnCdQKlq/cMclrHOaOa92yxcZxv6crQAuCqK5vp2zIn9VcFF30Tqi95fi
tpGSjwqm/uQai+7vlwN2Ll2uL0jj3L1zA8MjaUUgk0kTNFHnFDSS0LEn/XDipsmiokICb3+W3IVs
2AMlGJAk622WkKxoc6LfcXmZ7cxQ0/PzsXMDqlL7HkZ3JnmQHAoPI47LLs3+5tFGEfCq/tZHm4Ub
4x+gTWrn9s5EUnN4QsjNQcOgfzqAJIOCdpgdr7VkJe3UZbpIdzI2NDZ2lEfPuW4f22Mv3vfU6W0u
IuMBMf0GGWQJPLWJDoK3BB4x0RyC1zoXO5t8oc6llXN67dWyvxgQ+aKtwoBT/5pqPV11c5imUCEr
4igwEIPl726lb+lR3s4tjmeeFYfS+CPVweQ93IWTGXxb5aKzrSIL6McWGEGn2Sv6E9QZ1mcfHO1I
YvgTzeTFRVorV/EsSr+BvHJ+InI4RM2Y7dSoX1IjmZs+MUGkz1yhoDqR7qhah3BEJ7Lm+UdQm9yV
+xRrFteigU5+V6biBfFHvIIKC7/KCV1vfn+6Kr5biCI0/Heuq8lNVkvL+NbmFL06M+sNsxa3+akQ
JiDhEoKRTAjdK1mnkZboivWFtDfKIb6G5nIIy3CCJKhCwkLGpcdPUTwvXvqXuBoRzoBieOaOZuVz
EWCbcfpFJAPnUWyBsA4J34KNX6zjMyIfGocwGsuYTIdRW14DSVDYVn1FX+ArJQmsk+KCLd0g0Dot
EAs1uERsBRDKzMEujgmCecSOIpbvcAG85y6qmCWR/inUI4/ZepOyGCiMo9O8rV8DmNGHUhZkH66v
76kCJcWeWWrnKniY+izkGtLFEUWBGhRY2lTxCcyX4e1qyeL14vpiXO5Xh08vxdXVQF4U81euTCH5
McoY3Ei3IipbHE5nE+iEzbnQ4Pmt1Lai2YUaL9Qyrj7AZ9l/iKFFDlhvKE4BUdJCSXhRtNYfDDaE
w2u7u6D/Ud/CmDon0dvK9Vl8VM67u8L85qdO8ARn95hgodThmqukX0M2+NDFLFYTGDI1E6RReTOW
dVkNUIeFUzozbqYCKLmgQH0DuQSQYke6oxztCNWJDUYtH0ZZ08EvVb4mGLCWZq4lK1P/E+znM0rO
WLcSvEAZ121H65kAmfJfHKnomSiGF4xxAo//CPoDXxeVH7AL1xMWLxcTW+TYEd7LZKgQ2qkseq/o
7fW48h1teRHgGaz4x+z94y1GoPmZh3kOaMDQ+T+Pn296HcwMTt2rvOb8KiTvwJQhjtEIjFOgPGrm
ba7GkeEhZNflVqLf8BG9PgzrVvAkF8YVIiHDWDXRlhlPqwQzsvVlMmJoX0WKSmfLY1sMBYXWtffe
N1p5RShBL4mdckd0JVLBiBVFCTnUuf+KOofyaVgox9f367/tLCkBEyqNATNkqmfvoKb4zeolPp/7
VGAOFbbTRfR41QqcewnmvoQac8DvVKFVs0wsC8+3QPMkMuHiiCp+e+Z83D0/0GapkZB6BtWurG8x
+vaSoxSLQWP/lLmnKGIy4qWXi9DgYB47oAaOhRMuaObDR9yWtcALgoM9KnHvA/DJDyUGkKWORsBR
f5OG5Nv5MTMeTKFeH3RRYRd8XdWFQZb1pl7BnuNtFtvVW6vp9o/YRQvghxQyV0FQFqM27ib25SWc
yq3+jvVr16enpxRabEdrSyOjWOHWE0+dBiQMtAvSQbSoDPlunJVPk6uYKZ1uLQJuAZhLUo3P++iE
Qq3rvzD4bjNh3fxM7AZs7Cd3g8L5HLMa+FJ3ErxhMbf5wAGVs55OZgWbJE4qbsVAxtT3jUM1BNQm
DnpPgL896s+l4XQmQufKfF0JCpbr2W6228cIciWPg8XaFRwH8VSMTrSlzxsUvmFZcjihEk9iPvc3
VtS51LIK6nccR+7Td4HpebQYaM4v/pvmbJ0U3TMcma9dL4U6MVZyLFTPTvq8g/nqGHsU+NLn5Edh
+qZH5SYSsZgEtCYpnAhLKyich2c4ZxiB3sLaINZNoJkgfvtVf29VCZ3QGV4DZtQQu04cm++mMvbU
KvyC7mlS4In3aSKqSEoXck6+WnLvgvDWkVfFd8uUT7L7nGt97HM/wwVT08t4MN7+QW1iACW7xkDa
pGAIX7OkRP8ivLKh1MqAXjRBSJC31MhMkHOcnT84DngFo7kdHWSkEDjkbDJGzO8L+yCOKraMBFJJ
AdYzM+YoTE74sidNth9/dviFqYHOO3ipu+CjVbGJoHJCbiXItBihiYPTDM8r5bCbZc2tTl05U40V
kYlgBKROeBGYuLQJ7QQcocr9R+qSVyKxegZxQoK/PlOyutOP+YhL++wbx01jsFZ/22XnXR52y4fc
wCFsevVnRQZo1ezAOj2leVA8fCSjBTFDoiMIggCfa56MdhuqYfk+doSatj3lC3IEv07uwfEFQXQB
XX2gXZnfzcaUD/1vBZegp8/ZhDZ+9s53oEbFLtkxPvZ0zJJM7+4FLQgc6oy1q+yKSauvhnU2N8zV
ZrAaXhHo2q4VWvcMXmDqzUA9VSlhguztIx0kj/NzLF9ZvVwvAAjvKtKM/J59LllKR+6CtOW4Kr1a
GJACXYysZq5IHBDYIyB16i+GjaASE+fW5fp361i+Ynm9KvLI80ZVm7tsLnkVj3/JLkfkceY1PE1X
4Oq1fJPAfh0WFS4ba1l64GpdSHtEd3ldM1bLUN5H+SUP5Rky53Xh+30PXCSMsgo0Pm3a8ksminkU
kjsqIhdDeS72Yl6LipkhUCNWjk0hqL7u82f1PFIDFnVBZkJLJC+RtdAfyh5IPtRKd5GDUreN6vrH
24A/gCS1jWZrQLg0vt2R0Ah4JE0mmzYLJtk+UkBU1ijErfeDjajkVG9dgbBUA3DH41TZ9q9CDBZ9
ozyZ/2fXd2OMBD1EdGaOc5tWYC8RMhPb/vjSFzzdyaA8UBHjDj2kaQdom2M3SglVaLdyls3nZ63T
VPM0JdZE36r5ta+wO6qC1aiRphjJs/v+R9DNgIKAij+6ZMnFVEKiq7PKpA9UtT5Tkg3tTgkvGcVL
0mMb3fbL3SGnFZyKhaL+jePdmhfghArfZJFaNG3mrSZeIxtFBhK6KFlQqNUEJF9EhizIzHX+IlTr
ah4R1XqqxRpRfy1ZUN08Wkqzu/IG2vFaGpdZd3wunUoZdm9BFrANXeTuXKXgONZaJwilVv5+6z1n
qMwhQ0X+V2Iw+hngj0JWAnoOnTm9HWRTi6lgtTKOF1OD4H8NxvLcI53UcF3dVmE0jYvSi+CeusCf
o+d81Noic669OsiJY8CfY7vXm4+Q3XhgWNslII678dZ+cF8u53ccbJO+FdDZKT9LDbeZtf0X05Ok
1LZ7wjnYoaHot941Q6EkDFlqwoqLZ4cRTKYwU2zz/bwqaxR7jk3+zqR7jYhrZ2oePJAYzx8RFCeX
RjJaHHzp17gZILS6IcWnGvkStcYbG/HEbBu8akowDPUF22VQ0SuZF6fP1DJm9JhFNDNaC0rioN0k
ssJzu+VbKu6aBzHdapK/3ADsOx5syRUKUpZY2krLwuyIKZcpUvNCUk50aIzsDXB8bSAhl+HaYW+L
ubWxm1ywdyJ2s6bZKzqH553xiFnnPIdyG9bEz2E2FQKkuFykbQlHqc0omc6x7SLYvHLtO9MhtkWn
0zq4TRTO8GbpIPOntvQn1SNn8AP7UwpvznpGi5YM/HDhVGBes8aYZ7qUuF+FB9hEL59WnX7AluYz
q6IZsGhSH/YMiUSarOGyECOvPt23TyqEpCD+zbZ4vRrY6dP2rPJUnBJAV+m4d5IzkYGmbiY0GnOR
88CMCSN4AXmAW09kDzTG70tg5P+ulcENssqEbNlCRwDYKvJRhkTIvEWXQWS2VNPpaBxl86OHso1s
zglv7D/onG1AvuhfTGmfDNdXHJj9FJtDAQ4TkNrtdCF9GEAa3v1WqpXtleedju8F0MNpTeXdNRSL
2GX7YBCOV1JH+ZRp9/FIlfm96zexSjJC9cv+QDSGh0yCOOljt4xAG7ePSkj01qlLhqErxwTwa/zM
WV9QAscrQNbErHBal2Y8hCj1NVNVhtUzH4iimiv3ZG/zG6QvUdljaDEOrrL81XtNVJgJywMbDkkr
vmYqlE+Q/4YDxoK2D4fRgcDxpRZSugk5YmXfic36HKoNAmneTlKSSjJTpgS7/AB+jfEk26qY3D9y
tc//MgKBpVQ3LCB+ca+JIS4EkBaC1PIuCgQ/YqfhZr8qRhN1lvrnL/iSrkqxZ5XBGqzU7v8Cbzsd
5gojz3uUe8lZtKRRecVCbfwxA7/8tfhYMMLosZ4dTvi6XxvyLCa62J7CSB2dKa0rnOgL51fn5rC/
iuvUqmX7vAo5ZDf6V5Y2rRQWFtqJx2XoMZ576MTKZ37MLLTHiWosVcWFHE5yRdl7p/7MFJEzMEC0
qLqHIaGCaUsvOajgcWUHxr5HSD2uG2orSf4+fiOuGVDgwW3Kg2J2yKDGZ/m0EqRp1W4kqhVl0ne9
s2ipcT6bSK/FY8bvEA5c5PfqgSbcgmeglbTxWUciPl5V+4rLDgsVotScy/DQk9aU/HNExMPB7EcU
gxEVJV6sK1YTdToJ1qzayKXJrHBJEfpQ/Q/6pcJkbQTmbMOkyYZAYMLDq52XJi9ZpJWcdLhKvdru
P4lRHYQw7gdGfmYjdgSaNy1hD1+4GPVIVas3cSWxswlAkQsWEqmyY+ZNLfPrlxKGMrjryhIgpfoy
PuFH/hdyOLPeAmSDfAKC9krCaA/moZZ3qpzR7nVLvOLM78PZ1VUR/fLhX0SFrX7+kmAYvDGGMgxt
pOfhr3wyt8OGWjXWiEwq3AWUTyOxp6XbgTB9o22R6VxtnJFzEE3Y056SHs+65Ure2bKQ857V+t8H
rM+K6Ysv2CXY0dLYN0a50c9Brt/wBYwzcgXmeRCrapK3DboHvbx5xo7FC6La3c3mErmsmg5szOX/
n1IDqo3R6i/cYQXcZ2cG5sEu8ECOolt+kjVrMzndJJatOzSt3FcI13tZysIKVn9TAxE3mzaBB5l2
faIWkGXBjY76c6b4g4xOeC4NPrFWNdJiMLuMWOnlcnTdIRwcpHV7cQMK8Z7mAorpozq4JE677bB5
hIDi/TtMlQ3fCfI2wh/pbVM/dLIfytDMIHhKj/nBDiVgKUQFueKgLGkKOaak+STIT1DKswx8oUns
swh+VQ//s7ibZuy/WlmAHzQ1GBKqVbkoQRcA8Myx+ODl8K/k01medWjn5///BE9VAO1ly9u8hDB5
AK6Xy5VYo2EZ/LAoBnwW2U40EfaeqjNy6jKwWXQy0m1yHC2+/LUca3MSyEBHP3bEhxPD0GlFmcOq
TNqcqBM4pyTM/Vh5RchCkXDhHFZwSfRWanOtr0WGaTEHDum0HnL768DmJ6OwJZF8PH77f2URo1N7
rF4ur2CJElt0uEJMOkj0Fc83I98BK2BCRkDBZMIfmmOHNsEVntLpHGJ2iHWLMwHtj5DITZc6zZ2k
o3UsMXq+puTAZWEYtCU0oh4Yfju7SKGDRx3Vj6M6xzCpFyuMjZPtwatFij8yZ9voHxWmr1oYkspk
7bQgntqhH5u8AzhpFbXOOwm7yHuPPFiREnEy+l9gSdG0V7RzRdxA+pk2UqBYxJKbv10HHsAUbtn1
kPtfgLdFmnoINepzNXHvvfXqOzxbjLWTOf7T+PQetxLFrRPTH9pWkci/rLE2QdIXkfUcEuxFkgZQ
3m02F9AFYfs/BaQYp4W5pj34Yov3Qy1eW6UH+iaM7NWMlF6BSZUb2a5xvXHXUxqKbOD5L2wlGihE
ZTeW01OG9GwaB6UDUdPosFA7UkPff3gJVJX+ox1difvyX8NH07t6Ex0qR0Pyt6SVdpbE1Oj9J9Bo
PDweyaubMOPKpfP4kMtFi3n2nN2XOXGEbLPu15PiSoRs7+MMq8cmUILZVbqvLKt5bB1kLBadHk7s
hLRS/ksJtrDdj0DmvwIfCeBfFrQG/dbmOq77iErpd2VphrXHUmTt71T3Zc4lqDWzKTvmJbNPirLU
n8SAWoHr5wuLZtpIEpJzSdJ5vZ1S4qO1S30jXSFueotf+u9qXZTEjAtPp8V78pG9UddB+YkHjaah
Ml0utoQzlAvND3JRdQRPVrM233AhcRdlykaqVNWSMFxxDJ0wSEOAT8dOFrhexy+KzuyHvxyRuGVr
nhducecw/Uu7IqrFG0VNTQVkRH7T3sAyMleIxD9niTXcUg529QMn2asK7kIPGS3O1++A8UV3R8yT
Xy/U7ItaUXbu0vqYFWHFJyxNJzDgmBJcC9/jEQTaIroxesagpfRPW+OAKPo4hcFwL8PdOq4AMllJ
iE4XARq07cacysaPEmiuiBv2jY/e4Th+u349E2tD2HTT4xwC9tNIaIYt1EcpIEH+v49VjN7npj/2
Td/xGfkH6kwYP9+wwcxDkwJ/SOCJWg0oD+foI0H+W6BAjNuStSVXCO+njV/4rW6a0AfWkXRAPKmc
C+Dpf300osO6q+eTBGR7TKK+kK7MyZoRnNP6OqVFpIZEB238ZmM2CouKIIDZa8mBKPp/lQxGAHyL
yVo046LpLgUc60cDK7YDli6LhcixXAxEH0MnnJoG1jFzA35m6rR0fwke75JTque4umhiiPA8yZi3
Z4/9omSeD8NoxcwlB8uT7KC8W8euyoDel91cmrgX2yrNfOSLrLmyvCM6QWEAJWZWXaqbE81bZTvg
6Dcir6sZLL9eacBEYJkpuKC0HUVLu27bhPIApUek+IifXg70qYuaCciC1gWVtyyIwvKTRDP2XIe0
lUDYcPQnE3fPJttdtiOWjg6bpeGWaKrzQMrXsP9ynyuyRZ2yODT5wXYg2iPpmtplwyFvhnHGt5zG
RRb8HhOwSyDpyLXRTPytm3JvvCQ4vGPC41yx4JoPz6kaMoZnKDNceD+UPJgq9k99gDBXNVLjwKee
5lsCVI9/58nrbWtTecfK7iDQ4hm6cY1nmq1VqK/P/hWZ8jTFBm37eyGci2wktyxMmNt8VA6J+pVX
NE9ti5ectWT1KlC0WnVC+jkeblQlBed5Wvt2S8NrFK5T+83Fn6ClzOjIFTt4tNjxru5fCGRFNBJE
Oa1HFT9YKpPO1Fd85hLt+5yr6xeg6Xylzqh7vrzycWHkEAx3pWnSM38tN9OSLX8FCNL44HWb6IRA
GzhrBif7TtDEvSFZo3IydpGTCLAdS3ItqFmAjjWzUhMaf5k8Tfb4puLGDwjwwcZu+lzQkG3jxc4d
HyPXDKM7ujywPMrfYgphesTJLYHhrL86hE+ujgI1S5Wh8QaYndPWCn14QCnU9u1PnA7CHrJxnyDm
qJKmB73zw9wyGqPp8B6ne5LFd18knsTnV8GtDNiGgvE0kL23L1LMoMpFYNgo64AinFo4hy/20xx9
HTA4/NXN5AihhxUnYLXQocjPVLo7NxfXwrIrLHVMzZhVHF9c8btSmjRA06Z9ex290tNxE6apAKB+
mHktsnR1NUop+1x2tNW9ZBMjbQlmedJCG8nP2vYOGukOke4g8tE1h7GtB7L2f1nILqk8K/PLOpsS
e/yd8OtiNj4wmDP5fcjIQV5nZumnAb3QLvf8/t/jpC+HABLHz3ZvYzNT42napRpagodFTDRea/XU
nscSFMF0YdRln1wPoRBV12D45j9WpvYKG221agiEdI9UgrO8SeQgUux7NQzyrs0klUcbdb8lXRwo
xZ8mOOfEvt4MpInHp5Anf50L5JX9NsK5/r4olDFh+tBv+qTN28FnDTWHknl2nL5Rj4GUqoQ8wcwH
j1cqxXUy60OKZl3P/uesjQ3CuRuIGFuyo/afsY3BmIZxwpu5XOPxIhlSWJ469fFyl7rUXzT36vGC
Z4WskOw7qvLR5ZVC4chda9b8oIK6IuDUdWuqeNttEh67uEZ559oC+4oZmvUGInZlpRIIMd+HdDh4
RI0c8eJXkl7bNpwLf+Jnu3+tHgDrMEBM172X9Ce90/TG9WExjt6s3trHO6QJEWcswNgT5YbUVB9H
jCzvqqgg4J5FQ5Vf7oFnCTtLueVkQrUEkA+e0zWjBYtazqqggafuOVa+rHrWeQPDmOT5L9qCMpZ4
+3wgv0Rmj4rvCJwar5iF8LOvXRkI8Dxt1E8GP7Jie8hdLIwdO3TkwKp3dGVxDD4iCXVj3L7By7IB
E+lA5xkuJLAYjR1rYl6ShSre/ZyfFDXMeL+oKHedTEKOaWp+RWxj2jQYNCNJmXvC4yE2aoeuvvtS
ialPSP5w/2q2uB0PT5fImtdo9UnXQlR37tAW6kJOUXb5tlaE8ECHv5Hr8CdzWiV1kMz9J50JoHhP
5m5keWPSWZ1J0WXR8zafWr1V3K2OlrsQdBe03nCys6/DzoV1DPI9Bf1q/iupRNg57tgfdSpGVbna
l0tWVHCMee+NC/gop2ZJntOA08dnUK5Np5zFJgJcM6lLstFvp2tieAXgDVzvu71QEgMiwrXQUo7J
7J2jjP8BNCcVYgQs6/JpxiRZdXM9gJHn0g/KS0W+iuh9K4aJG6Vcn5cWuOptEl4TEYrL1QeI8YHh
oIWbW75sWbnbmc3Fv5AOcigF4OqL43apAOQKTB7USNs/v7o6stjssGiOPHrImZ6TnxfYZwI8rj7A
3wo85Q6Hk9ab5Kwjaqfup1Rj4BAb39gqdZTJA/fKaa6j7ik2qtTYujz8hqP1zmeo0GS/EZeSFJsY
Gfbjf28QM4jt5dddidlmGmINSbeju0JMhyBIPQhioa2DAnXajorXBt6YKHsYpXpoMFF0p1PPmjvg
gW78QulAgsF4TCR/WyyxBxlsn3jLIYHnbcAUkC1bTy7wcpQeGGJWB09YAsmFuXe0zE7lO1qAVpLA
xzqQjUasVjhAYjM32L1Cu7EaNnnPyZKCxyob/FQm4I7BpCkclqdIH8psNWigjA66FKsLb2FdCK/i
LZx1iPBBd6NHSrAMSTdPblLoGY//RDQnWrEdLWc0JPWtZsBeWMpZ7P8k6ozZ0Wz/ZCyEwTfyl1Du
XmfcxtNx+KvPDWauv5lbhn0RYtH0mV9+doubglnL7+TS0DJ+EbZ2WpWLfajfJw9xvbLKUK6OGWS5
Qz/NkCjWhvxtOMHI60Xyr2pnxNJ1LwPatW/B0FO/nXn74MtsCOTYL1LV1Gmq0CjrzUHJU3um8QbR
ZqnKsvXrXPa3WU85bajP6SxhEw54SbEQm18l9zoUTIxMMw/Ky2vsf0OF9sxgk0mCXXCx7YtANUQh
SBOmKcBfZgRzju6NciBJlaaz+ha0F//LiWR2tNAvBJIf37mORaAcjqJc8iXpr5tB9UmQCeuZp0lc
VEhcWuuYn9hfQ85quJC0PyH+NPTGioxk57NdFjp/BpIwHpHc8l9lGLe7j4Yo3VTQOaRq/X3F4esI
yUS+AznA1+Wmi2leC8o+pYK9l8bHEwVIYxYFnGp4h47Uer/XBXYDsxBNiIpTkCmWmOtZksTYmE87
HjtYikraH1yYvs4nbfna0bnwSX2JCSVHpQIkeAWKeDDbHJTgnva0z03XyY+h73ia/0xtw0T0yi90
3JGOzMLFMTCaroRJ/BzKhNAMe5Kx2qwb8TDunNwB7rKCylYfXa6fJh0tEr38KzOza52B2OU2MhMI
qDZRZpSDlzbNbci0KZAJPlyotjpB+ZvyBSHJKiTABR/XfU5H4DVuUiFbzG1jniFIJ2kXhLTFVANQ
XOxooyrMV9l2fboqvozJBflmA26pCNE5ZR7Wm1uqsIeFxebQHedhDJzxMij4W3QgQww9FZ5ld5LT
UeBRbFTRFpD/YImIH5IilCVFK2eYF1pKcEPqLi3+fev1zWV6MR1vFYKtz2GWPaLnqkaoZpUFon5d
kdd0Ww43R8hLuNn5U51yAWWM70xz6t3lT13Z2Ws1roarV6mbHC+jJLmPKkONxUJE/X1rscGQ23oC
Tdu+7ksiCsxPpySF7T9zZ8BMrFZh40dqI0jokiX40HayXh9+5hUD5cbAoB5imeHkJi7f6bUNeKLN
luhhPENZ/Hj25HSotUj19wb0aSbFDri/P0fPnjK68AxpobNGk5U48F55dZe/JnCcke83AYM+xBHy
irzsA//aZMXWiUCS8QLSXWWWTye9LeX14Opx7y8uO9+f3JNQHiCGEzpLDYy6q7wLWVMMRmkndPU+
oBRasxPPDorCXcMPNEVQloapMpuh82OM42Xk62/spa66sXqDq4U0u7F+q/G2D5N2dMLLcaC7ylXy
uoHEBsHwHwY4aAwpqj1t/E+X1p+bMmmRfufK3+Kv8YxsxKwFHYE0uqjx1+zWAwl1DuxsTJ4IRLUT
4a3WydlWbsjxifOM/SPmh4Tlr/j0cPugp7m7WKf6m+XLXPPMS2R75Tq0al3gn/8LTI7wNW1AYI8w
qt3Y8N6zh2S+f83s/IVV4vKnde/yiLJcthygdHTbtaCvd9+/OByvHOBDYMnlyAgiKjS9ZOr+ovuZ
SfaZxb5Af+F0fxFtWCsOQXo+V2jO0hvLdzR2mpyEAMFTjMZSO3DtwjUUaec7QOj6t0AdisalEjln
Sldo22M/Hg6/2T6aufhEmdwdnCbbuVAIUjBv2Ep/MclJvhEaS4k/0192KzwaRaz6KA6FJp+nZsEw
QmDWILURwQ7x0sMy6a3AgE6IlL2+sKdQkREa+JqFAXoMn6TTGY6sMMP+uJ/U/uz9I6B6l7kFpISs
DWoWSxPSt+M9K6Qy2oKpJ7Auu3vMupsUFIsz/p8zyYi9oXbS4WackCzsAXwdULFcfH60OcwIqog2
+9twperFyAh++50Sq4U5AR41XKa3bZC0xAuJ74KtEyrsBSZyLDR8Koaj6gU48RpPBinLRpo+JsMM
rv8nFiZGD2Pdm9KWUHPXqTehU3wqBCFoOlrMdLCJmGEOTeryCU83TwnsMSyAAA+XTOOpKdEnpSvL
hMo465Hzdor5BMsvsDc1BkcfPxHjEt+i4Xh0OSQRhKpCpmza9NXnsqNETfvbnb1DkVbuSd/KerQL
zKJoAgvemHjO38Qw9KQsMWk7TZZTzD40ltV8euc8VVjLQ3/wqr4GsXklUV7yF+SaP53knlJ3kYon
3r5BzWQ/wmh7EMjibHLpWSBLtuYAFSwmgwBU/Zj4yHEPmR9QY9056zq1YiLvU2axIaJ0AoBqFctc
NuedT9E0gvx+V7gxb8VpDEaLamgVeDp4A/rC4dCrVwjkTvMcsTswuC2QJwWm/4A71fuOBFhWtctI
t8odTc0xq+EDawkhitZRMJl8ty57VOAF44E2WgTd3hMonp+1YZ85eofVi8zi51N/Z3tTb8gZ4wD0
IGiuyFfocQIH8n9G3KO/qQeePvXd9wp1sUCdIqLryGBKGPFBJ6Iidn2naz2Et/hvtVkgImW5fAz4
4+c6phu+ZZw2cLllujm0UuQNhayC5xxPiA1f0ew39nl1z17soEyErkUIFvnQCgMdvt5OZ0SJ4WpU
2v+E28jvmbuJnoi7dQwEmyhPtqcUdrHPQPYgxmop0AmStse7kXXtHYssGNGwkWNLwVkJzELXrYbJ
0ZC5gMZdKEU9/EUcEx1qgHCZV1pHULatqabTam13yJc87U+4AV7j9rKiTd3MDNbLKte+87wGb7F3
ZBbKsJxqfyk0S+1Q8qY71+ITJwGdVoQorICC5AMMg2G6cwcppNLX9Pw1QatkA+NcXgHeqh7IfKNo
W5VFZmtX4uSEQn5V4WU9znoq9wBtuIVwq/c4u2yI8K/oIV78If3frNCz79JeDGmEYXs0jvOT9o84
wNoHSquA0cHHJFxqcWiZRLDIzI1UosbeMp2beHxRgrmTS+Ag90KM99sfrCViAkoDlVp9H/YIA1Tc
6gGZr0NZae2wB9MJLJBeeqskc4TL6T2bAgO9i/nEX25qTHIOC5HaqFp5W1P5U7WeezdJCPkfA1kz
/dgICYSEZzS2dm4zwAdwg1QPyOeHuIhEifCI3ZK0OgCM5226xXpUiw4gGO6Stb/ItoCmcSgHFkr9
/AA+8wrn+5rYhpgLCJVlkD1DpwlbnHU1T1UKR1RaQBB9QeTWIbw95QHHK/uzsBdmHGuY1MQNE1Qs
IjaNlEYgTzHrXezRF8OBRPwSdERtMX6yjCrGUvHhiuaZryG0bcxQJJrhtr2oPgZS1wgmEx5JGkQ4
x2RgNKAu9TJXWBlD8gikF0OFHizglfNY16AF/lqoPINZNz/yF2aFJwtGYDQYIoM95vxf7AqGbM4L
eOQXAe2sv365oPF7R8knTGqgdNqIpqjUL01vC2mQK95POmOBo5zqz41yH60ZLzw2fNslgFbF0JH0
dOYd6hsuM7Yv9IBGzsooxf+VyEPfCcDZ56molmBF0PnNgpn7WkmgrfHNjmrLpJ2HLOT+BK6yioZe
skL3HO0I3ro3WZO5Waz2Wj7UJmx/0yphfFRc7Q/P/Jzad30+N6F9sPVUVrOf//P7CrLdPymReCEd
bkz3y6/QV9oD+rObVXldQmbbG2OUZPuKxind9SkqOn47fh3eLphuGpalQBkn+HT2Z7K3KSImb6l5
i9KEt1oco32pRAm/jLubfi6WX/9VTX6E+e6sZlP2rPUWDKihaJ6MnUTJZmy6uMuqXZZR4Z+G0nCk
affT4aAKvQ83lblQxpGtLrn+ir2jKzSk6SQLRwnvEpsGKspRhzunAoQZ3FE8ev7+gUOhWjVkmpHO
7fhkE5OJYrHT/CGUPQoe00fST9PuWMvcqmO7cAWCammbOHN1Od1WPSD9P/oUptBlo0ehkjoG1Taz
Btm+/WGynOcz0an12XQAJSG6pUDT88e8meZZl2NmIuortbezgQ3Xjfiq1NOnkzpcVjESHnSyc6d5
5F3lmOhQx3JYKuJGsKIbSXX/JUiXtpfDbbFlUiGWuvP3TSXhxZyBL+KmiYm3Q4PdfJKH70DKRsBR
6VB2Mp9EmhuQZhgTcR3FTAwB+jV8f3zcditULSpl2hJ7iPWreHoJHU8m3XT2iLTDt5YdNLAdpvHr
f29sKS6+tGoT7dFRF+4sSXSJlVOBukeOo4dZRlDCqVpxw8t48K5Gz5TWUDNaCDX+r/l/NsCin7yZ
jk+157bTtPqQipqHQBuo1VyIkSqPc8mzXg1p/BjztrZ+o5KZNSlG837CnHYXyTzzHAf9aF4KJ23T
tT+Dcin9KyIDTwFfPwcymXFhwOaY0BYqqbL0Gzj25a7r3eP5xqr75DRpL8PGSLgy1FeyVMrkJbDJ
5GpX7rgMe5f1JMM98kqPWFOrNaFwMat+w4nJhIBNkr46QRo4MRAiuwDqdPcy8EHlMMt9nGsJ9XEm
V8d6cqubONmcx+7zMqeeaT3tsQzJJ43IQpJot800idCZjbB5q4XQxLzF+G5Rk0Hj6DPq5kwtX0oq
E/iSAraNC2EJRNgu+TcIUH1LX6EQGhdm2eUAg2WTW3GAWoeqQHgvAXvJy4o0xScEpQsyN3om5L4G
n7jpVthPUoFUgqI87lYCH4oUWXMATgl4+zEwLz5D/n3gc3ICcqnP9s1sPVS4kpF0AwlsRd8YGiu8
zQAfVyQ4wWxrpPakN2fpkMKXmHfiydChK6nsrf8gefF07l35btf056Z//7FCP0wcFSp/oELlXxvM
Fgvhi6ckB1tWW/WaMibAKwfqCr5o/kJ1kOHMXKQQB+amt2HGALqnqFGN058DdvmUtr9nv5vh2HSY
DjleoTVsaMl+lqOdm4uIIFqZub8GV26uK2JfZtKf4J6MVtUnZFdH9eFys4ZnIKhPsM6gUfGxIDHK
S6sxC1hpFeKY0D/CilxTZVdIF3dBUBPSsjEKVKp2mkBX+9+DvZ01/4Nku7Zzcx/w9iOgW8rMNK1A
qhlHABB2AwIJsAFAHKhqxntvo7rb9+Ko/fcYKpkyLq1t7rcEQfBqshqHV7vudqbxd890CSarZudZ
AmD72GDE2m2V8ojNj3YTCK/7Rn7l3kTXSOX81/jJh/GCfxtJcopNJm+sKScoR5Tal7RngFRu8Yka
mqdCxH9xjr50otirH3jvsx4QfelijxwMFR1csVtiaFoGBK01HTzsJ+Bz/Ez/sxsGfljAkj+RtpQi
iKZ3pARF3j0ZTvPuE0LM0qjBo3JQvSi1S1fCMyn8DmUVYNA++LOuK0qSsQSP7cJE+pPLr+d6+2qB
3GYiA04V514C+p8UjSfbsn4728ywbCCgBRBO/DrlVaLmR3bUlabsEJ8VooIvIFFUGF5Z7YDy/JWW
VW6b3MTqzbYR5UjvTI8k50DIs0TFrU4tEAdmSbjarNSt+T+gcVYA60DpTAW67Wx+mt3aRbNFTuf7
CWcJxySZNYpBb3FiiNqu92yXQ0x90/dTc77ssyclsAj/RpiebmuzyCSgmC0QOeS16rUQ+7osNvcE
0NERf16p2k0UBr4Z595lKYGk071vy5UPhNW/v3I4OSHKcBZY5y7a5+uAFyTrM6CZVjYQCtE2W5Om
QEF46o4A5WcAPcAl4SfJvseDtEjHxkUmvdqbQZH0PcorF13LS8xOMfoQz/GVSV0ubLi7/LR4RSqo
HQk1Fa90Y+J1d40uUd2YlcjYuQ8i/PdMMBIybQmeVJsB2LYsDxktMIAN0xbmRT+oHDVrOMM75C0X
dptu6m/ck6S1YMrWVFk0cqk3oolOtsEcTGVCXnq3kShWiondYX+5OlrxqFGAvVZuJLaCTUGod3bk
m6swRG9kflRN/a/07+sQVnKAf3frH5JhPU+NMB/Pplo9C7JCTbfS2EgeunIaKieSbsLB46ge1tCC
LP21SLxw+wngc+efYdtqJ8IAAJVMotuwp7OalJI2HcvDBg9wwvERYpcoZKjbt3ygPScyx1cBMOiw
wvLmD9tBzm1GhVPDPIq5HHRKl2WhPS/LHeZgQ7rJ9T/eMbkomYto/4eni/0O8WcxUlvX9uWVNzWW
YCRPxZ8CZowQbq+rGeNtXh2rRZ5StpWPI1fUDNW8/JczPD3tdyTdM403zWKZ4NyA+IgZJwbiE9LS
Tz6mWxc/ETSrV7HK/W7EDreVSMIda/xh1vtinxVzBcPwrJB7v7u96r++8OFqSoGc5vkn5tXaxFQp
z0eFi6SRwfPThmuBCBxAZLbSxRyZ7XCzUfd4WjhTz6QDDS9VfQPWiSjhvvdbLYF+jxBwI4NuXIH9
URbuwjWZFD7Xxb6JPs1N3IaRe2o4uXBOjEkrftbchm2Gt48HNzc/im+NY5EhwvE4dMvQUazqo2xI
9uWbDfGSjPZZ62/EuSDYY5oA2+GKlN7bt+nrvy2tw5X9Y1ufe1ZvrGYAP0QUUijCHcTVHoLxWmiz
xbnFqO67a6Q524QCm9iYeWwUtbyAHyfqq8vINByhbMpecEZkBPyBTwEvRtlECL6FTN2b4DKxXNda
DZmAZoiJrf2qIFrRGEZny026JPp3clQzXNtr7DLNDBzEHKQKLNWhJLG1c4aZ5fgA4DtGvvslcEnp
ht8jP9bC9p/N/Ln6z1eRQRs65j7cf+XVIVGIXtiTmEijGfp7qYQAHVG8rVvvv2G0RbWlmCkIP6hr
hhcaAEhtEZ9lowIpn/Ni+ERu7t0z+LbucBnLzcB3S31iHKxZQw9+2MeSsVh9XNiQfJLjQB0IlRU6
dpVwgMbff/N0oA5plZA2MNwEU2DPStjfsIrOxxbJbijYF6pjLWazxz/beT6oVPgaiU10AUI6iocU
4GiiCiztZD5uatUsaakJhcDUNT7/OZUEuxkf0y+qFhpffm+fLHV8UXErXh1IoWazinA18rNZpJQn
OTZn0wwqf8S3Z/a1O5rMBBLIAYRGLQGdpee0aPOFQagdvOjy7zbcl5qAy4mOkwjb9aiUA0KA2FfH
C7JEbgOOQMAx9uDKOH2a1fLpiKB7HgFdrIu/AMo2GeGjOufpNTZ/6dxZk138B+k+iXmM+byebTsX
wpFCoXfhT2iLYlTmGfxCJ/QhJXReCxEz9YfFkoH3sNqahF21DlgrRR152py1E83xyc9GkkT3bkky
V5HUpKdN7BCLrHY5LbPEFyaoevzW4OeUaSLTeBW8wMXP/Ba79aqIWxwA1W6St/c8nvhOtZX6b3Y9
VKvEhjJgeC0Q+qm8ZnhXftZzCVGXunuDhimkQBF1CQyXotOSGNPUcnWlxnawHEj7XlPQ4eBca8y1
DTuNaeSNsLj1xcwNbKSRZA/+jNPaMZ5u3xWvaqOGrYkcLhvCiwCqG3ygDk2ss3UzhVdx1WFA7V9I
roe5IdWr5CxjpQmAIEy5aR3095CTgpc5OIj0B7ujM3+YU+70WCwbliQdHxfehD29V/gIsuR6pSie
v+g3IJrmnTW6xK1Ov8j3IRyLGW+BBJtU9Ae2PEIoSMNV45QP4ZbTgk9uWnj2oI1vFlsM7KMGxd1X
JWSHXyHT3gqbDH6SHstwZRtaYT0NHWCA+2mydVmJFWqLsAP26tETF3C0PtH9DcZvlt5rFdiByxgY
Ct6uh6wsCbX+/9oOaanIAKa4y5wHaQ/uovgDcTFh3MBt9bAFNITRp8LK2SmmHR4kSkCWTYO0rovS
oF12VaBGcuODV183HVurADFSluOymNWTeHcKjcgK/TdPiUjB0VLOcOCQcbJejyB35Wp9feGrahmy
EzNb0QWe33rLwpAQ0LzyXB2bwHMxyY73dwsQZKHFOeE6J68EX6JaTe3AcTdzvQcGfGViN2i5W8ca
k/tEQ589K9v3dCRYQIjwTTSoaxL439SATX6gI067FZgFP7h7FfpvAkMDCSwzdFaS8dSxiweYdxlL
YN0GQ7RykXrfeib84SFxX9mMDeDaWDdz08lYfEIa+8xbVcAlvDM4QCo5pZvqh/789zizR9JWeLRn
1OP7YdgVVZJpi5HkU/wuzZoiwotaJlo1Af5MpW9PvEVEClElbuacFFf4wsMJdHqXfhPZBM0+2ftB
DzmEW6f//+nQS7OMBL0lsgfWlJvRxhBl4JrG9BhRTyH3nRIRuHlAQjgw0C1aQfVgwE0L6DTUbREh
p0fZx1ZPNFb5R5KFmHywGMmT1Lp4fATRgiV2ttkGXPtdmFpsIk+is7jCCZvkgwi7+6LSLM9rMD+o
RDCbjrdarsA+xnqOwyhYfAEPZWdtUJCbu/LmMRBf6V+RjXL2CP68gbDDFhP34kU0xvtv43CbcJTi
uKiCK6I5lfAqDbULFg2I6scy0utCJxJrLGRw+4sOkAI3mAVlZtfn7Z9DhQpNZ+7iCDH703QWYTqt
Eh2TYI+XGMURR2iCgbxLNlEP1rgJlFk1aJ9tBdEgsWuu6KzDqCk6QC5WIMTWZ7QXS1s2awVdE/Og
UsBqedraLlkkpr3Eegfh4K5vzbrb8+Efuu/vhUYkFIx6jpCay8UyjsufoOp24l3g2mfiqfPez9hN
0tCLOGJKvZH4ABgx7hkZwromFCD31wfM+i+NtFehNNMDtmJRLd/uywaHzcAHWZMl4W/lyGckXOrN
3fgh8dXuqjHtpL5MgmyQOkyFxwpQSm9HNwZv4egMds3adCbyQIM6PFwtyaVn+W5IcmrS4JrFyF/w
1MWMDbNrk4ukLezgCGK8uLt8wbByj/h4njFPj5934n3aeKCh2LDdTMx4gwAF+iNcH1qygY0sCuT4
KQggkZIGt2sHm6IaUP8a7YxkHdgAVzVUt93WXDl6iaYezjutsXbX2YjLf/hO4bXvMDuzOTmVchSZ
7EW73eYXvNcaIM5HtcYzPq5h0W9iAK2AfVA+klehVVLzfwjvd15BOAwOj8/FjejfIqcVYH9xPiNw
AL8B07XRgMZvnJvtQHkgxPTfRTDqmZ8UBBzoVuQp36COaA/OsDqoDPpfQ4R8W4S+0+rBj5w29TI8
zwPfL0IIxX1tRn+gASqPdnzfSQOhiGXMNS5srWGi+SkZ/k/hju5Iy97nlk4Vyw90weZ5a1yClYc8
Ep5qm352m5i67nXNfU2zn1dWt3Db1q7+JXfCVfSLplo9UlPaBGpRQRqB7YezmmMULlpVwRZj3Hqs
xUqtR9mrv/zKA5uY+TWB6Hg2u5SughW2/CnHNavHpjrtQkhTvBV1EwCuEe8hWMwKv+MVr4+AoP87
rh6q19DBJKJauUuX4P/7etX5oTKZBrSpB2Y//dxMMCpaUsyuXxb7X4izQGjMI2GoDPuU88FI8qY0
k2o25PuLF0+LTIapHRIQSRUQ7GPTYI+hTKeNMl4ParqBf6xhvfdxDtsVE/w+YImz9LE4G+3bNsNR
b2yn+lesM1dDkNrBgYeB/vlgoqVS33wBISZqPjNT16AcubMRgQujyljNZrAm28FURvZHtbFo6g+8
G4thqS7Yj4r1zQ/SDqD2TRHvZAgL7QcRd5A7LxSqJB2uHRnDk2y1TiDDIfZflVUKCl5C7rrwp6It
WRJcLbU7Sc40cXY181U7wuQJJ6kh/N+8g1jdFq+L3w+9VYqGqxfQad5P1WeQ4hEk0oBkj6OCfD8W
KIykWVndjMr0dGAIMrg6gDFC6nqejIM6kq6EqEq+qtPs9FLqYS/Rblji6ORKwW9jLGVEHENsFNze
wyrniS5b2XWGQl+z4Qt2KYRXsuc3SY1gjwAlz/BWL9JksobmaJCaaUu5oOqXGgis6Ethh/+GuOW6
lcNTuYiOS/qnpdkYhu7608kyzWuvh6mqSeeVaaEXyDviqnBjaSovOuDF5u/WZrixxq9Ea79qcCzO
UyvRZbWiUip73Y0vKUpzL78kNIYhDVVF4LzWSfRi/eKuUcpuevcyV5V4NSe8MvbG4bWEJeyzI+xo
fF1yArvuMGtCJmufSc3OpOsGiihQMLXG6lrH/+4+jtElTP/2q+/d07umyFttE3LdS3f+4huyfsRV
oL4t7u8T7DZvTkIVUhxBbGlHbH/rVUE/i5W/HtXBfK/A1L4i8pLkam3z78F+5Z0vpN7ucm/8LkJ2
WRlHQ3/j5ggxyEW68YzfuKqsOv5wOkduLmCpHnJzebIzRb/0S8cT4WHwDwDloZOIO8Lp70pC4ALy
ONptSuSmOmHSJPaNW3/DFvPYS4YQf/r8UDRv/EHjFdFNXeaQ7tTlViA5IRSIZAUB8lqM2hXoxsjr
qSYHAIRMwE02THjxzhAMtSaFWvCnm2H2WkALgVGcssDd0DjUuUM0+ThyIr6ccnFAxjvLoXNCTiTH
FPxwqdvcWwSraefgv/xtxYsGlsncWnqryrqJguI87YKkIxmQJOgL/xo9wfVvvBRLkGJQGqI9AYEa
A0j6hrY/LmvSXKpKHkrG8E1Ofpa3ea3gttYePKSIO2TiB0np43lngsFrylKaK/SP9PnJZ8XYXXV6
o4USnhaVlXWJxU2XJYsXBSKgC0Vcl5gv+niBsSMkcA78/TB7YbWWhTrxLY2U6qONb9RmXTsTr9lb
6MIJ6O1Bnn5F7DWHxRqlYTEZjxrpzzsiE5FY3Qwb1Z+Ixj6Nc+aHdGPovqqc7xa2UPUk/52olMP+
O211xha/+ECIUom/vK7hD8QXiu8vtO8PuhFEHaJaJdlv5xPPIzryd2XzbH//nWMLgL/J2pKy0CA2
ElGhMt1WRlTHeV73CuMmJGEWb7cQwJKyjX1DWgcklMhamavyD+I1rAYniY9ECk430UBOO7Pb4XPU
W3GmZG7OdwroRTAJ8osGNBvxjDTZPjDXKxT993uzvGwivElHcI9pmope+gRb5rKJaeJCnqtzQsoj
xrBs2xL1Q5JR/nKNqECChhOsyLkcgN6c085+VwjcGcA1iTaN8eBZBkWCvy+160mgF/fKbFm2y7FY
X3wCf07kqAy7PwJx3WpNFZf0z9GQ7ES18kcLdon3bmWbMAajfo+gASEuC4L1D5A1j6lJ1f7OSkg/
HNxW12CNhDGsdtZL6fp3aeZab3VJ4gVQBUwVHKl+Gnus5Wv5JXdbyQrWdp6PtW5Q+08v3YXUDPct
BGLzkbSN4ZNzVaIJWDWxMCOsjDbhr9xg7oXApU8YMhn2GcUOrbz03/OCv5QgW6SfamZ+WaHqYOn9
z6LGSHZhh6AOK/o9c1W1+WzOvHtKf+oW0RvsLgCsiOO8ER2SNggqYEnJd4y13n+0ybMCEt8IUwDW
7qKrdVFy+hGCSpnHspXB+Rl6maHhunJSZ8Tt6/2RcLWhDxP06nBSckdDlvdEWVJ98WjFnXSQs9Ak
pAu67zY/yCcqMR0BtrecfNAcfD1Hnmn+pGluCV4LdZzBRE23B6+cdeNvFoa21XMXNdY7oCKOyKPk
RirSzpiPa3Y5HwYZ+8MZTdeSGxgdaWKBsG80PNeiHVHzcJk6kl0q5QCXVSArqBhfNbG4iHherON+
tcZO8CGhOF+LIbCxKSwsofVpsys1U/0vXLzx2eB8mZeFR27+ZRVX7pKlVo//K2hlrQyZGJYjqWek
We5A2Vv4CVQJRtos/FrhILRaQUfF6x4XxQUmOJMMVaJIDErOOvpYA0p+EDred2GfwSKFSy7NrOyk
EejESPB7BbIA5nOFF1Dip6jnsT2AN59pRgQyS6OqfY4DvoRB420RhsyXmjJhDmwfMbIoCZ1NDFWf
6JzeaMwXmNMUAD4YNHKx2eC/y1sXYrrZAd8UDSwf9FNDGR0PjyX6J20T6laHj6UnW4kp6ylCy4V1
8ne5jyFMKO22aJRZu4gOsfUgv1+Q1e7X6BGPohYGJETqVlcem4ZX55kTVn/lo7jbsSigZKbNNH0k
5kcro5y8voh/pTSj7y/3ZexvsBFi2Qph8UgH11QCKdG9GSp+nSYS5qB/ZqWW58yjNHSkzZaInkPp
3j1dxKUSqbSwnTOlpna0SJwOPX/RzVhXZpwh8nqd7d2uy7HLz9GropCfvjlJKvoPpDza4N2jIMLr
88gHdsP57cEMPCfIKLIFEyFcp+sDHYQlULq8K+8bS6QZJqTNEZiYSDRXEpQ4RIVxaqJszwvpfHle
gHDN4ykoBq0VSxALqyMJ1uj6K03/7I9+afZv5Hu1bDPGRaxe8a7ogHZyQLy+WaTXvYxFG1/pB7i2
88CQEpNkqOhMQ06L7BQvHIFdKG05OGeCwBnSh5M4lnWM6fOJKmsnZO4JgZFAddyZNEoc+5wN1g8S
G/bUW2h1qSNTdyDpPG+OU7qdT3ATTSJSvS6A1Va+KCkWtC0nZMnDV4Z8UU+FqUf5AqW/7w8a91wA
gv0cVyT+66E9muHgSdLnYLDKNIea920CMeu4vAWl5TxBllaITMTSJEwmIASl33xAxXX1PHxhSjeB
8Jgk0XOk8MV8Ir99LFDb0lrDkQah+SP0BJesmGpE3MpBeXS0Tm5Dl68i42FtiVVCEOvvXLd+IY4W
PsZpcq+QIdEyz0PysYPcRBYOdbw8CiRyYP9yHYuvIAugPxm9GbCnEl+l+y+JoN2oVNzjODngU8GC
62vrjIxKhvxTckXLH38eapKpYBezqtO9DiWp7KcqqyCP1gxNeAfkpJWhjGSRXsi0ndkN+G/e/CwF
qozyAXotP1KILWizMoakGEVnb2VDMH18+5+SSmkMz+7q8Fyxv5tjqxiaPp8G8PiYkz+YpNh4T2Ki
4xQwfNmyWh/PE9aNCKUx2iJk6zaX7N6sxT7R5DNFHhbr2GIiRzMzEINdMR1r6djPw7OmhVXoQPhT
i5bEp7pCr9VxAYOxQ3Ptgs3TdOKCIxh9Y5xaFhjZiorGX0BvHtFTOkVtYFPfvzTCwOrg2nNP5rCF
1KSbcJJjMt0Wbq1mhbHK/9kIedsiOx+s8ZQeC1rZbWr+nFl3zO9/9M3n7VhQxcUkW+FuKb905ETt
/qUS4fsRcc97oGdn/D4+J1uAbPrmZ9xfzqujP1zlDngcgh8iqJpdi04/GknxmTjsF4wJLZ+EsJyX
vU0HqznlzedNa6pYJE7A8ZCQ2zFWFLzfPZpEXjAFMMeRWOwrTwejvCXaoSoe7f0kzhI3eTC0+42a
jc7UECLTYcJBirEIex7odBMCAfPsyEClBgfuORES+LY7DfCEIvBhe6137lcGTXBVLlhsR4VWV//R
byGy2QgLLFZNbrQxeAxOZSCC0N9pGD+V8St20FJvRyx7VBB4WMx8L/IkY5IeMM9q4dgUzULXLbt1
vNZyc96+sBdxmk9B+m2FzT81V/Cs7s//n+vMBLnCh3vpqRYYouMQrBDeyqBbkl8gMTXkOkZVP9hr
qB1BMlGWfi/UTP7SyvbSI29klSvzwQfqacQuL5Lv3GOCTWyCHRB5YNAPKmiSz0x+X525y2uauF2f
NMxDvJO1QNvbm4134oX1obpV+jelhs+aL7BCKVEXbxgWEi2ytNDnDY6a393LXHEdf8tA6Pk1fYW4
zSfLLw/3xLEwhF5JaM/9Uzei1kMZ7Rmxdu+uauILFiDRKkNvR1/LC0/8RQy/AnjaEmQLIb8LYB9Q
q2jIrzlI7z00RzAsgX+KHswMbFlD6X4X3cppzJfFdPdVbZ6rvqmDIzb3yPTKUY9e/ND1ptBQHGHS
/5Xp0sIqyVfHoLU/V6RDLhY504iNVqoiMDgo0yLh+vz/tW5+1gqdRohsMzil85xkiexcycbmD2FG
w+aVci4Xu1EW/oAk4GN+nknkmXXkg6Ml1I7erKlT3O6f0g9W//oQR+/c/FrfyKEamoqacWLpHn/M
6Wef/8UfC4KysnbZVy0XLlas/0lXPLEix4kmT8AxImIyH57fv8tDqi6x+KefDP23sz6Pn7H6tE36
GBLQxYtfUk0kf537G85K+gnd2HZqrwEO3m9hdIIaOUslS+htxKVf9B7Pr8yl3EMk9EEOEodF2oVD
vevwsx9KZc5eU48EHk8nLQwde3bzcIgL59sv5iceoMBq0paecMwfrMV2sM0coYxriH+B+xZOeowN
ErscMYYH9ShftjzaeGqy2q5E5VoB++n8usc2n/M3ZhIPdo5ygIlNgrC/+JLLk59d49Tfx9JDULXv
9YR/z6I2BGIDv5bWGXPStJQdnfMjFPE8kmVjRTAl7xRgROUxY+OmKgr5klrcn3P9ei15yVXldw3p
3uo92m+cBC3/d3VHdbZ00QRfW9fJrP4K9IrbmkwNBSq0GExDVGcjSiEJDP82kqhdQJkJMJaUAE9t
k80c9cbi1unZpkjYf8FszWJQXTZL+2o3brhGMrNTQin0PK3tR++v4XH4GViWFIp/w6GqqdCwLhU2
qfa+nK/hMSFy0dlWGNTcolV5yzOzx+HULPyEIKq+Q1dl8MUBNzCZNcn3aQ8FC4aPeFDJ/Jq+AwLC
kg8UuXfP82eBPDklukEgYVIPZzfmCcbQ5PmzA5Z+v0ZM6MgjQGmCZHIIL99nttimJHUNMvAVCAvy
JvuWqzDJf2mCmnF7IhllNyPqPT0jXAirSqgHFUEraySc9YuRnKGE7EXkp2T58rQZkwAXS02tw3hX
68bW0m1xfYBSUCCyYqaWwve6RCWlXW4ztX817fjDHtT0YoUGzL72S2i5/DGRXj8i3qswNfaYh1tJ
qIXKV2sVlnO+/13TohvwFboWxdBQkzQ9UEZOWGk2Yl6aPqp8cnFxuGE0h5Ohv/gWRcgJgku0dlat
YttlMhy9Npfjxs6vogsaGThNdNVXg4ZsrQ32RstKY23II/Ug+Fhx/7D2af0Nz+ojPTwJwL4nl9pW
+RcpRbK6okiyk0NpuwCkzTkukcrtI10v5S4KbfoHI4bGYI7x1Pa75zhLSge0o8N1xyyb5ErLssvB
p2D0HzdrXZQQ6+9hM7StfXCKvX4PeJ3x6Ri4dT5I9vBjBN6jboa3voML9hbEgpDC9gU3TTxQQtZj
B3GC67j1o6mNlovMp0XGTMSdJWYgPdZmZp56WeTENxdMZzY+1/0cy6v+n6VhIYmleQwA0ql2jdZ/
CM/oNSHFFHSej9bFMjVGihur/omUkO8HI8Rd2xaWbaIDmHYCnP5ejk6ZLYaYPotJAkigBu4vO9jr
GkuuvnOk7Wh+x+VxBdxcownIxqXf4GBU3pZDq1LrCsYWkW7gvdVKQswBgtkJ7O6Xd72vZel/CDy8
jys6FpX4ZVcRTFbL0cKQNl7A9lgzOIUfwnIjutkJ13mk/5RANZdsIvC9GH62M5mMF+1ihhAbXOE0
v8g4uuOtvon9UrVDFdcnUUByqiAa+O38hz+OsiZR8/NV1ZhVKuaLO38+DbE4Jpj1Ns9RbTm5F5XK
WFVmWsHP6YBEQSOnQKxLV7d/U49Qi8HSBg5jTF3OzvOoMZ1WEE1qV626/L474J6aSAorygjxvIM4
yxJHUcNmrxPSfcIzSIqEuVdrWY5HyRUn7zO9sucIcoqnrlHlP8nELK07sYU8DR85ijXZNzwKRXrB
MDx1xvlkG5z3cRCrqOA2VbLWRXidycj9dblS3+hhZ1kbWvYu0O8OWgJab9yVZjOT/dHpQehwfhRx
otPUE2fSh0W5PJVafQ2n+IhQP1Nn+1Vs2P7zWZpH0Wubr4lxp+KomM3HjLykzyHnSwTN/r2DlbjH
O+IwGqNCZh0jPwRjGpj7gmsFitrEWw9tUwIJaN9uJwtQ4pxDFVL94mJnoqNADli9ox45GO2ocQBo
xMsKmgkCTt29uGF6uUxIw+NeyADa6rM46lne4d3yPfh2Wwgp72ph1J4VwMFyf7PahO3bxySIQODO
9mqK+w5easJzmzzaHvx5+LYJ2jrSlvO8cNy8V7i0ZcJ6hBuqWEKTxDaVOMbZd1WxAkg6V/CoIEsv
MCda4mnPSpNt1LGy9M61CadXgtOVUnMdMBn+QwxiaVYNSKupnP39wg7MFvklMwHYQlwG0ybpzF5G
urpLsh/CCGrK+RceAqrl/vZ17dhOG6L/tdnQYRCpM0mVCTsQu9jGEZHF+J+1MQTwxpT8s6qTB0bz
j9llPWeyAcFnkGXnTvFgd4NxnMc550kQrj5fsErRUoZKIK2mhCZ85lZLellRC15xcPeg7+cYFGeD
ToWTw7/4b2YKe6qloXa883bug7jAGzxqVxSiBSf005VFhrK+xPc9ABFAAZCXQLf5dRhjPa4xuptr
kDbPhXv3hXOXhT6MqpxjbmKqXn1lxE7PCzjXfrrQJ8lvLtEzsYtIf13TrHPyf7wRD3SQ5nKSfZp8
1heXQsey3e5oRStnZ2iDstDt2RjeOlffEgBReE/b1SoYz6h+mxLnIa782tPqSaxqO9efBpYFFLxG
Vtb6Cplk1sdjwhwC5HcySsm+RMArjz57XUWmW3+N6i7cy1gGUQXrxxs+kQOQP3cCl5XHWneX6oiy
tLSJa1W1IXIvZi/G2kATuBRdldt3azOsVlJ7bHaTCHqQxtJX/gw/TgvG91YDjboxBKjSORTpWe/A
DetJ4H25G/OPospXynX/G8pEz4DhCUQjqbOI8ax1tqOvockl81CQTzKmRNmsiwrXQ752I+sa8uBu
y3QIhSMl3jeAjdbytB/DwvDdCWizS8FReHK4inCWP9uh48IPeJtdXtxvZURvndwTQTG2oCDcyQUP
NSqMPFFtaOCu6z7jr0G3fxtxc1/wWrnCzt8I5+xhovMd9TONsw1cJNt9mYIBTUjamhkrEFBcanHO
vU+tCUobFMEK7oPCW+NwvI2tqfoXlbz0R6jQlAd2JPO9BCSyh4uOfHR9CHH5aKZx79RQEBeG8jE/
W5Yq87wCSlPg9wdpVt9mM3GtBNfxrMUbd6c3oK9OU43yWNYbGAym76Tj71WCnHMVSWHj8VlTLAXq
VnJ3DTG4w7/tPJ7f6Dck+7GHb8HYRgy+l2qQ3L0Mc+JNB/JkEFXYocpZORMnGOxRmjGt+m6f0U4q
ycPrOHQGosM8qeYxNDVeJ8unzraXVqPqDKDGU93NU9dPevZ9mEbZa84iEhyxeorNiy7/Iw+qVJjy
yshGmq9QaSf8dlHOzvdv2B6+D4+1eizIx3YuietQSqNqgVrQwPi6W6KAM7MG82HEhIylmFmX2NEy
JTq7OndQ8CxyXTMIcmI4WoKeAPJVuKOAFXKpqM5ua69k8pR6KJJc2jZv74fVThh4/haE4q1resky
eqKdWExYQNlEFP6TVn99Cyw+rjggH5zGIlGtfa14N646iCDRYxU3EnmpkRLFV48tN6Nn4aikt2Pn
49jWb0torZSguhVu5Z0xIELE8bS/Ljx/HvyypvmfQu46nZRWDT/CAHPxToBRhrfHT5CeOLa4Hg9y
cwwLeh1v3ngFu6m19Q2yvuf21DfQjpRyf7yKubrhvj+ZrpxCXh2YgwuLnVpi6GpSl917pau3/qXr
6feMjhLZmYwYkyCwBV94DTVmK/83iE4QAZyv8rUQVwmD3w7AwHtjJbSs+5v2PrQ4NVZmBHyHDpZb
qMs5QRBY+bGWPsO12GxdavAGompo37TleXzoa75bahBZpESwCK7n2atIRAzKDi/WcteIzkw6V+s4
RP7R2Da5DqJ7aKg1VB0JSD6RvLopCKleF9kdFXBIuHrPE5iASmZuMD/0EN1ZLOjow7sNZ0dlxXCM
1fM6HAi+PhpTq0Kaw49u8dScZosn9A1xPkVf9JkOEoan95v88G5nONTeLIrFPS3EZoCV787O8Rv7
Dl+qVnCoGVoW4NKRulAv0CqFA8+wBfXsTfWanCaX5MCIBsTAKgPLvdZ/7jv9Ken46zkeQUaowcnH
A/hwD33LKo7QgV+y5/xEBbhzouXNQnkMSZt8lb5+slyPd9Lt+cWTI9qcGyemf5lvlufpYsTgyI9N
O6WI7YLKMKJuU2atxPDDOg+WWsbNp9hd/P6HLHqEpOX+Phzi3eHwWuEeuumCRyH398fEnEUw5bUP
WKgvzuolCX4UO5Ed80LHu015FDDHBDu4j6ZlAhEr60F25jhXMCzyY82DBYP8u1hzWqa+jpiGugRF
DlI7eieU+84CQBJHRdPWBMdwOqvbkSCaRItC+nMpHPT3UeUL4gjuwJsSq8RhBir2B408uI7RFDbI
LuqHoxcbSBz9Ty5fU61cDuL3FZxHhtJTtfs49TKZswFzpivOjfjTOOdnzuZkG64Va46NrH36epIO
Es9n7j5E7swi9v6ibC/aXkhX6aFNP0wYgUPWDpuDGx9/C6JpmUNcSs9uVtB6Yung0hlqu70Vh00h
mJAamScEnz30mmTz0sgkOZ5UHEOs4TUEpADHLdux8BIzyAN04O+qvAB750dqGvdqOs04M3p2fGlE
Tut5AJJNTty3SmoYiD6afrirp6G/8tHOjzXPTpn/J6rnC0No+nlRQrA7gnAkwvTAAQoKvi2bfqbD
hRZmfV7ci23CbyRNxNMqsdYCB2AGzEBJi/51Sp6lOaiRoBPHHrloY0XUmfmnh28fsui1bfdZpa+S
nYYeK1ss2ARuqnikCJHMg/n4y1knoncQrSNF6rg5D8Njc2mjHef89mO750gHgdB02BPog54iUMLK
3/5hvJCsZ121ubMHn7eju/0/8mMl4iIoXp4Y9ZNjLj2bcMMuvKYfqRtjvBB81yj6klo3HyxHdeR/
80LrZwUlu04SC/k07tMOVzciK7XR67bX44WntARtDC6sFVlDpuYncS5+cIIOaRZF8TM4rkN0TwQ+
M9b6HBivAlzkJrUa+tek0XDks8JcfaYRBJ6264Vo6XZSQV4G5Fy4QYOqgNEU45LwwKRwUbOUri5h
p+3TWYrQ1D/BTt63hv3tezyvGlU2PamjuBjjwoVIJ+EJGS5H58Y07kMBYDnnNXGj7wuTOquOXNk8
1WGkQBWs1HT3+RLhIfFwFhf2P+Y4V/P1RcjdwnCUxvdsHrHc5R4kjRM7K2bI3F/eI38cKXtoQZXu
Uq/VrCfccTMupu2gFpMI3ZXXobOeykU4FzvXpC1JqudadFPxqd5NcVSUEGA5OCzB52YIbeI8f8QH
61YByT1Zls2SG16pyvhWbGsrCyHH/jnmYseALnccZU7oDhAtYXUaYWbTf0LFVDhXlkbi3cMPJIOs
JwgpFXJDda4rXZ0hYCYYW4H7egXLCK8NXLfXpKpGzwI0m2ULoCPUEXN2oO4V5FLxa0PQklOAwc13
dI//rSCx90hJX5r3nuzafjpLuD9P57Gcxd2utABN3idMjBb38tWQSeQ8L0B2QWsDWOZuwk6+3cEC
cP7MbK4iCpcOkkVQksv6udLl0nsL33sAjz3OsQeH3ZakLc3di4SxcEhywP2Tu2isy2XG7EAjmwJM
9DKMwq8DpsPruFy4iyQhABwh0D6HbnBM11gQ8L4yvatOV7duEHGYZAOZ5AUeMrZiaoavth77O9mb
w3ujU/sHupSnXQTsdU6/xgRtT4z9Zt/z/aAfsYJybMPSG/mMYAE4+NxgTi8DzBGaOcUQ7GsAA00h
SMktwBdNS2VOlX6WNF6zpNXrzLdkPJ3uZppH/CnEaSQCfHy8Rku6AEpHUSDpyeSuVDona46Tv3Vs
MYncbdYdy0R/HRw4H76MXdP/tms/hsYynpNU3WoJhbR8O7STB/q+lMoHFXmdJpAgbDjMFesSxmfS
kQd6pqDvdvYboPnu3nbFroHZ8MTFuIWzx68x6QuV2YZJJZdorPyR6cDzrEZSfbTWpN7B1V+t3oK8
5IC4Y0FNaHNS+V4dmkTSsbgFr7uCcOUIQQv73BKRPpvcro4L1L/IznOk4rt7MJ7McD5nRcG5z7TU
qePJhFqhzEZjQJf/93KTtUji9vX8k6jgARatKRnyNjjhw/PLiwp1tiysxk9w8jbGRA4FUDoE2w51
RHX7nySvv4xMbfksxoU7ERJq8olLqUKyL+a7kBaR
`pragma protect end_protected
 