//Setting the arch of correlation

`define def_IMAGE_W      128    //the width of input image
`define def_IMAGE_H      120    //the height of input image
`define def_CP           4      //the calculation parallelism of channel dimension
`define def_DP           40     //the calculation parallelism of disparity dimension
`define def_IC           32     //the input channel number
`define def_ID_BW        4      //the data width of AXI_ID
