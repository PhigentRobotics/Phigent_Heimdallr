//=========================
// Engineer:  Wu Di
// Email: 
// Create Date: 
// Module Name: 
// Project Name: 
// Description: 
//=========================
         


//AXI4 parameter
`define def_AXI_DATA_W                    128
`define def_AXI_ADDR_W                    32
`define def_AXI_STRB_W                    `def_AXI_DATA_W/8
`define def_AXI_LEN_W                     8
`define def_AXI_ID_W                      8
`define def_AXI_AWRLOCK_W                 2

//AXI-Lite parameter
`define def_AXIL_DATA_W                   32
`define def_AXIL_ADDR_W                   12
`define def_AXIL_STRB_W                   `def_AXIL_DATA_W/8